magic
tech sky130A
magscale 1 2
timestamp 1647362286
<< obsli1 >>
rect 1104 2159 198812 177361
<< obsm1 >>
rect 198 1096 199718 177392
<< metal2 >>
rect 1214 179200 1270 180000
rect 3698 179200 3754 180000
rect 6274 179200 6330 180000
rect 8850 179200 8906 180000
rect 11426 179200 11482 180000
rect 14002 179200 14058 180000
rect 16578 179200 16634 180000
rect 19154 179200 19210 180000
rect 21638 179200 21694 180000
rect 24214 179200 24270 180000
rect 26790 179200 26846 180000
rect 29366 179200 29422 180000
rect 31942 179200 31998 180000
rect 34518 179200 34574 180000
rect 37094 179200 37150 180000
rect 39670 179200 39726 180000
rect 42154 179200 42210 180000
rect 44730 179200 44786 180000
rect 47306 179200 47362 180000
rect 49882 179200 49938 180000
rect 52458 179200 52514 180000
rect 55034 179200 55090 180000
rect 57610 179200 57666 180000
rect 60186 179200 60242 180000
rect 62670 179200 62726 180000
rect 65246 179200 65302 180000
rect 67822 179200 67878 180000
rect 70398 179200 70454 180000
rect 72974 179200 73030 180000
rect 75550 179200 75606 180000
rect 78126 179200 78182 180000
rect 80702 179200 80758 180000
rect 83186 179200 83242 180000
rect 85762 179200 85818 180000
rect 88338 179200 88394 180000
rect 90914 179200 90970 180000
rect 93490 179200 93546 180000
rect 96066 179200 96122 180000
rect 98642 179200 98698 180000
rect 101218 179200 101274 180000
rect 103702 179200 103758 180000
rect 106278 179200 106334 180000
rect 108854 179200 108910 180000
rect 111430 179200 111486 180000
rect 114006 179200 114062 180000
rect 116582 179200 116638 180000
rect 119158 179200 119214 180000
rect 121642 179200 121698 180000
rect 124218 179200 124274 180000
rect 126794 179200 126850 180000
rect 129370 179200 129426 180000
rect 131946 179200 132002 180000
rect 134522 179200 134578 180000
rect 137098 179200 137154 180000
rect 139674 179200 139730 180000
rect 142158 179200 142214 180000
rect 144734 179200 144790 180000
rect 147310 179200 147366 180000
rect 149886 179200 149942 180000
rect 152462 179200 152518 180000
rect 155038 179200 155094 180000
rect 157614 179200 157670 180000
rect 160190 179200 160246 180000
rect 162674 179200 162730 180000
rect 165250 179200 165306 180000
rect 167826 179200 167882 180000
rect 170402 179200 170458 180000
rect 172978 179200 173034 180000
rect 175554 179200 175610 180000
rect 178130 179200 178186 180000
rect 180706 179200 180762 180000
rect 183190 179200 183246 180000
rect 185766 179200 185822 180000
rect 188342 179200 188398 180000
rect 190918 179200 190974 180000
rect 193494 179200 193550 180000
rect 196070 179200 196126 180000
rect 198646 179200 198702 180000
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22834 0 22890 800
rect 23386 0 23442 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24858 0 24914 800
rect 25410 0 25466 800
rect 25962 0 26018 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29550 0 29606 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31114 0 31170 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32586 0 32642 800
rect 33138 0 33194 800
rect 33690 0 33746 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35714 0 35770 800
rect 36266 0 36322 800
rect 36726 0 36782 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38290 0 38346 800
rect 38842 0 38898 800
rect 39302 0 39358 800
rect 39854 0 39910 800
rect 40406 0 40462 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44454 0 44510 800
rect 45006 0 45062 800
rect 45558 0 45614 800
rect 46018 0 46074 800
rect 46570 0 46626 800
rect 47030 0 47086 800
rect 47582 0 47638 800
rect 48134 0 48190 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53286 0 53342 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55310 0 55366 800
rect 55862 0 55918 800
rect 56322 0 56378 800
rect 56874 0 56930 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58438 0 58494 800
rect 58898 0 58954 800
rect 59450 0 59506 800
rect 59910 0 59966 800
rect 60462 0 60518 800
rect 61014 0 61070 800
rect 61474 0 61530 800
rect 62026 0 62082 800
rect 62486 0 62542 800
rect 63038 0 63094 800
rect 63590 0 63646 800
rect 64050 0 64106 800
rect 64602 0 64658 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66626 0 66682 800
rect 67178 0 67234 800
rect 67730 0 67786 800
rect 68190 0 68246 800
rect 68742 0 68798 800
rect 69202 0 69258 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70766 0 70822 800
rect 71318 0 71374 800
rect 71778 0 71834 800
rect 72330 0 72386 800
rect 72882 0 72938 800
rect 73342 0 73398 800
rect 73894 0 73950 800
rect 74354 0 74410 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76470 0 76526 800
rect 76930 0 76986 800
rect 77482 0 77538 800
rect 78034 0 78090 800
rect 78494 0 78550 800
rect 79046 0 79102 800
rect 79506 0 79562 800
rect 80058 0 80114 800
rect 80610 0 80666 800
rect 81070 0 81126 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83186 0 83242 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85762 0 85818 800
rect 86222 0 86278 800
rect 86774 0 86830 800
rect 87234 0 87290 800
rect 87786 0 87842 800
rect 88338 0 88394 800
rect 88798 0 88854 800
rect 89350 0 89406 800
rect 89810 0 89866 800
rect 90362 0 90418 800
rect 90914 0 90970 800
rect 91374 0 91430 800
rect 91926 0 91982 800
rect 92386 0 92442 800
rect 92938 0 92994 800
rect 93490 0 93546 800
rect 93950 0 94006 800
rect 94502 0 94558 800
rect 94962 0 95018 800
rect 95514 0 95570 800
rect 96066 0 96122 800
rect 96526 0 96582 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 98090 0 98146 800
rect 98642 0 98698 800
rect 99102 0 99158 800
rect 99654 0 99710 800
rect 100206 0 100262 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101678 0 101734 800
rect 102230 0 102286 800
rect 102782 0 102838 800
rect 103242 0 103298 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105358 0 105414 800
rect 105818 0 105874 800
rect 106370 0 106426 800
rect 106830 0 106886 800
rect 107382 0 107438 800
rect 107934 0 107990 800
rect 108394 0 108450 800
rect 108946 0 109002 800
rect 109406 0 109462 800
rect 109958 0 110014 800
rect 110510 0 110566 800
rect 110970 0 111026 800
rect 111522 0 111578 800
rect 111982 0 112038 800
rect 112534 0 112590 800
rect 113086 0 113142 800
rect 113546 0 113602 800
rect 114098 0 114154 800
rect 114558 0 114614 800
rect 115110 0 115166 800
rect 115662 0 115718 800
rect 116122 0 116178 800
rect 116674 0 116730 800
rect 117134 0 117190 800
rect 117686 0 117742 800
rect 118238 0 118294 800
rect 118698 0 118754 800
rect 119250 0 119306 800
rect 119710 0 119766 800
rect 120262 0 120318 800
rect 120814 0 120870 800
rect 121274 0 121330 800
rect 121826 0 121882 800
rect 122286 0 122342 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125966 0 126022 800
rect 126426 0 126482 800
rect 126978 0 127034 800
rect 127438 0 127494 800
rect 127990 0 128046 800
rect 128542 0 128598 800
rect 129002 0 129058 800
rect 129554 0 129610 800
rect 130014 0 130070 800
rect 130566 0 130622 800
rect 131118 0 131174 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133694 0 133750 800
rect 134154 0 134210 800
rect 134706 0 134762 800
rect 135258 0 135314 800
rect 135718 0 135774 800
rect 136270 0 136326 800
rect 136730 0 136786 800
rect 137282 0 137338 800
rect 137834 0 137890 800
rect 138294 0 138350 800
rect 138846 0 138902 800
rect 139306 0 139362 800
rect 139858 0 139914 800
rect 140410 0 140466 800
rect 140870 0 140926 800
rect 141422 0 141478 800
rect 141882 0 141938 800
rect 142434 0 142490 800
rect 142986 0 143042 800
rect 143446 0 143502 800
rect 143998 0 144054 800
rect 144458 0 144514 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146022 0 146078 800
rect 146574 0 146630 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148138 0 148194 800
rect 148598 0 148654 800
rect 149150 0 149206 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150714 0 150770 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152186 0 152242 800
rect 152738 0 152794 800
rect 153290 0 153346 800
rect 153750 0 153806 800
rect 154302 0 154358 800
rect 154762 0 154818 800
rect 155314 0 155370 800
rect 155866 0 155922 800
rect 156326 0 156382 800
rect 156878 0 156934 800
rect 157338 0 157394 800
rect 157890 0 157946 800
rect 158442 0 158498 800
rect 158902 0 158958 800
rect 159454 0 159510 800
rect 159914 0 159970 800
rect 160466 0 160522 800
rect 161018 0 161074 800
rect 161478 0 161534 800
rect 162030 0 162086 800
rect 162490 0 162546 800
rect 163042 0 163098 800
rect 163594 0 163650 800
rect 164054 0 164110 800
rect 164606 0 164662 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166170 0 166226 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167734 0 167790 800
rect 168194 0 168250 800
rect 168746 0 168802 800
rect 169206 0 169262 800
rect 169758 0 169814 800
rect 170310 0 170366 800
rect 170770 0 170826 800
rect 171322 0 171378 800
rect 171782 0 171838 800
rect 172334 0 172390 800
rect 172886 0 172942 800
rect 173346 0 173402 800
rect 173898 0 173954 800
rect 174358 0 174414 800
rect 174910 0 174966 800
rect 175462 0 175518 800
rect 175922 0 175978 800
rect 176474 0 176530 800
rect 176934 0 176990 800
rect 177486 0 177542 800
rect 178038 0 178094 800
rect 178498 0 178554 800
rect 179050 0 179106 800
rect 179510 0 179566 800
rect 180062 0 180118 800
rect 180614 0 180670 800
rect 181074 0 181130 800
rect 181626 0 181682 800
rect 182086 0 182142 800
rect 182638 0 182694 800
rect 183190 0 183246 800
rect 183650 0 183706 800
rect 184202 0 184258 800
rect 184662 0 184718 800
rect 185214 0 185270 800
rect 185766 0 185822 800
rect 186226 0 186282 800
rect 186778 0 186834 800
rect 187238 0 187294 800
rect 187790 0 187846 800
rect 188342 0 188398 800
rect 188802 0 188858 800
rect 189354 0 189410 800
rect 189814 0 189870 800
rect 190366 0 190422 800
rect 190918 0 190974 800
rect 191378 0 191434 800
rect 191930 0 191986 800
rect 192390 0 192446 800
rect 192942 0 192998 800
rect 193494 0 193550 800
rect 193954 0 194010 800
rect 194506 0 194562 800
rect 194966 0 195022 800
rect 195518 0 195574 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 197082 0 197138 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198646 0 198702 800
rect 199106 0 199162 800
rect 199658 0 199714 800
<< obsm2 >>
rect 204 179144 1158 179330
rect 1326 179144 3642 179330
rect 3810 179144 6218 179330
rect 6386 179144 8794 179330
rect 8962 179144 11370 179330
rect 11538 179144 13946 179330
rect 14114 179144 16522 179330
rect 16690 179144 19098 179330
rect 19266 179144 21582 179330
rect 21750 179144 24158 179330
rect 24326 179144 26734 179330
rect 26902 179144 29310 179330
rect 29478 179144 31886 179330
rect 32054 179144 34462 179330
rect 34630 179144 37038 179330
rect 37206 179144 39614 179330
rect 39782 179144 42098 179330
rect 42266 179144 44674 179330
rect 44842 179144 47250 179330
rect 47418 179144 49826 179330
rect 49994 179144 52402 179330
rect 52570 179144 54978 179330
rect 55146 179144 57554 179330
rect 57722 179144 60130 179330
rect 60298 179144 62614 179330
rect 62782 179144 65190 179330
rect 65358 179144 67766 179330
rect 67934 179144 70342 179330
rect 70510 179144 72918 179330
rect 73086 179144 75494 179330
rect 75662 179144 78070 179330
rect 78238 179144 80646 179330
rect 80814 179144 83130 179330
rect 83298 179144 85706 179330
rect 85874 179144 88282 179330
rect 88450 179144 90858 179330
rect 91026 179144 93434 179330
rect 93602 179144 96010 179330
rect 96178 179144 98586 179330
rect 98754 179144 101162 179330
rect 101330 179144 103646 179330
rect 103814 179144 106222 179330
rect 106390 179144 108798 179330
rect 108966 179144 111374 179330
rect 111542 179144 113950 179330
rect 114118 179144 116526 179330
rect 116694 179144 119102 179330
rect 119270 179144 121586 179330
rect 121754 179144 124162 179330
rect 124330 179144 126738 179330
rect 126906 179144 129314 179330
rect 129482 179144 131890 179330
rect 132058 179144 134466 179330
rect 134634 179144 137042 179330
rect 137210 179144 139618 179330
rect 139786 179144 142102 179330
rect 142270 179144 144678 179330
rect 144846 179144 147254 179330
rect 147422 179144 149830 179330
rect 149998 179144 152406 179330
rect 152574 179144 154982 179330
rect 155150 179144 157558 179330
rect 157726 179144 160134 179330
rect 160302 179144 162618 179330
rect 162786 179144 165194 179330
rect 165362 179144 167770 179330
rect 167938 179144 170346 179330
rect 170514 179144 172922 179330
rect 173090 179144 175498 179330
rect 175666 179144 178074 179330
rect 178242 179144 180650 179330
rect 180818 179144 183134 179330
rect 183302 179144 185710 179330
rect 185878 179144 188286 179330
rect 188454 179144 190862 179330
rect 191030 179144 193438 179330
rect 193606 179144 196014 179330
rect 196182 179144 198590 179330
rect 198758 179144 199712 179330
rect 204 856 199712 179144
rect 314 734 606 856
rect 774 734 1158 856
rect 1326 734 1618 856
rect 1786 734 2170 856
rect 2338 734 2722 856
rect 2890 734 3182 856
rect 3350 734 3734 856
rect 3902 734 4194 856
rect 4362 734 4746 856
rect 4914 734 5298 856
rect 5466 734 5758 856
rect 5926 734 6310 856
rect 6478 734 6770 856
rect 6938 734 7322 856
rect 7490 734 7874 856
rect 8042 734 8334 856
rect 8502 734 8886 856
rect 9054 734 9346 856
rect 9514 734 9898 856
rect 10066 734 10450 856
rect 10618 734 10910 856
rect 11078 734 11462 856
rect 11630 734 11922 856
rect 12090 734 12474 856
rect 12642 734 13026 856
rect 13194 734 13486 856
rect 13654 734 14038 856
rect 14206 734 14498 856
rect 14666 734 15050 856
rect 15218 734 15602 856
rect 15770 734 16062 856
rect 16230 734 16614 856
rect 16782 734 17074 856
rect 17242 734 17626 856
rect 17794 734 18178 856
rect 18346 734 18638 856
rect 18806 734 19190 856
rect 19358 734 19650 856
rect 19818 734 20202 856
rect 20370 734 20754 856
rect 20922 734 21214 856
rect 21382 734 21766 856
rect 21934 734 22226 856
rect 22394 734 22778 856
rect 22946 734 23330 856
rect 23498 734 23790 856
rect 23958 734 24342 856
rect 24510 734 24802 856
rect 24970 734 25354 856
rect 25522 734 25906 856
rect 26074 734 26366 856
rect 26534 734 26918 856
rect 27086 734 27378 856
rect 27546 734 27930 856
rect 28098 734 28482 856
rect 28650 734 28942 856
rect 29110 734 29494 856
rect 29662 734 29954 856
rect 30122 734 30506 856
rect 30674 734 31058 856
rect 31226 734 31518 856
rect 31686 734 32070 856
rect 32238 734 32530 856
rect 32698 734 33082 856
rect 33250 734 33634 856
rect 33802 734 34094 856
rect 34262 734 34646 856
rect 34814 734 35198 856
rect 35366 734 35658 856
rect 35826 734 36210 856
rect 36378 734 36670 856
rect 36838 734 37222 856
rect 37390 734 37774 856
rect 37942 734 38234 856
rect 38402 734 38786 856
rect 38954 734 39246 856
rect 39414 734 39798 856
rect 39966 734 40350 856
rect 40518 734 40810 856
rect 40978 734 41362 856
rect 41530 734 41822 856
rect 41990 734 42374 856
rect 42542 734 42926 856
rect 43094 734 43386 856
rect 43554 734 43938 856
rect 44106 734 44398 856
rect 44566 734 44950 856
rect 45118 734 45502 856
rect 45670 734 45962 856
rect 46130 734 46514 856
rect 46682 734 46974 856
rect 47142 734 47526 856
rect 47694 734 48078 856
rect 48246 734 48538 856
rect 48706 734 49090 856
rect 49258 734 49550 856
rect 49718 734 50102 856
rect 50270 734 50654 856
rect 50822 734 51114 856
rect 51282 734 51666 856
rect 51834 734 52126 856
rect 52294 734 52678 856
rect 52846 734 53230 856
rect 53398 734 53690 856
rect 53858 734 54242 856
rect 54410 734 54702 856
rect 54870 734 55254 856
rect 55422 734 55806 856
rect 55974 734 56266 856
rect 56434 734 56818 856
rect 56986 734 57278 856
rect 57446 734 57830 856
rect 57998 734 58382 856
rect 58550 734 58842 856
rect 59010 734 59394 856
rect 59562 734 59854 856
rect 60022 734 60406 856
rect 60574 734 60958 856
rect 61126 734 61418 856
rect 61586 734 61970 856
rect 62138 734 62430 856
rect 62598 734 62982 856
rect 63150 734 63534 856
rect 63702 734 63994 856
rect 64162 734 64546 856
rect 64714 734 65006 856
rect 65174 734 65558 856
rect 65726 734 66110 856
rect 66278 734 66570 856
rect 66738 734 67122 856
rect 67290 734 67674 856
rect 67842 734 68134 856
rect 68302 734 68686 856
rect 68854 734 69146 856
rect 69314 734 69698 856
rect 69866 734 70250 856
rect 70418 734 70710 856
rect 70878 734 71262 856
rect 71430 734 71722 856
rect 71890 734 72274 856
rect 72442 734 72826 856
rect 72994 734 73286 856
rect 73454 734 73838 856
rect 74006 734 74298 856
rect 74466 734 74850 856
rect 75018 734 75402 856
rect 75570 734 75862 856
rect 76030 734 76414 856
rect 76582 734 76874 856
rect 77042 734 77426 856
rect 77594 734 77978 856
rect 78146 734 78438 856
rect 78606 734 78990 856
rect 79158 734 79450 856
rect 79618 734 80002 856
rect 80170 734 80554 856
rect 80722 734 81014 856
rect 81182 734 81566 856
rect 81734 734 82026 856
rect 82194 734 82578 856
rect 82746 734 83130 856
rect 83298 734 83590 856
rect 83758 734 84142 856
rect 84310 734 84602 856
rect 84770 734 85154 856
rect 85322 734 85706 856
rect 85874 734 86166 856
rect 86334 734 86718 856
rect 86886 734 87178 856
rect 87346 734 87730 856
rect 87898 734 88282 856
rect 88450 734 88742 856
rect 88910 734 89294 856
rect 89462 734 89754 856
rect 89922 734 90306 856
rect 90474 734 90858 856
rect 91026 734 91318 856
rect 91486 734 91870 856
rect 92038 734 92330 856
rect 92498 734 92882 856
rect 93050 734 93434 856
rect 93602 734 93894 856
rect 94062 734 94446 856
rect 94614 734 94906 856
rect 95074 734 95458 856
rect 95626 734 96010 856
rect 96178 734 96470 856
rect 96638 734 97022 856
rect 97190 734 97482 856
rect 97650 734 98034 856
rect 98202 734 98586 856
rect 98754 734 99046 856
rect 99214 734 99598 856
rect 99766 734 100150 856
rect 100318 734 100610 856
rect 100778 734 101162 856
rect 101330 734 101622 856
rect 101790 734 102174 856
rect 102342 734 102726 856
rect 102894 734 103186 856
rect 103354 734 103738 856
rect 103906 734 104198 856
rect 104366 734 104750 856
rect 104918 734 105302 856
rect 105470 734 105762 856
rect 105930 734 106314 856
rect 106482 734 106774 856
rect 106942 734 107326 856
rect 107494 734 107878 856
rect 108046 734 108338 856
rect 108506 734 108890 856
rect 109058 734 109350 856
rect 109518 734 109902 856
rect 110070 734 110454 856
rect 110622 734 110914 856
rect 111082 734 111466 856
rect 111634 734 111926 856
rect 112094 734 112478 856
rect 112646 734 113030 856
rect 113198 734 113490 856
rect 113658 734 114042 856
rect 114210 734 114502 856
rect 114670 734 115054 856
rect 115222 734 115606 856
rect 115774 734 116066 856
rect 116234 734 116618 856
rect 116786 734 117078 856
rect 117246 734 117630 856
rect 117798 734 118182 856
rect 118350 734 118642 856
rect 118810 734 119194 856
rect 119362 734 119654 856
rect 119822 734 120206 856
rect 120374 734 120758 856
rect 120926 734 121218 856
rect 121386 734 121770 856
rect 121938 734 122230 856
rect 122398 734 122782 856
rect 122950 734 123334 856
rect 123502 734 123794 856
rect 123962 734 124346 856
rect 124514 734 124806 856
rect 124974 734 125358 856
rect 125526 734 125910 856
rect 126078 734 126370 856
rect 126538 734 126922 856
rect 127090 734 127382 856
rect 127550 734 127934 856
rect 128102 734 128486 856
rect 128654 734 128946 856
rect 129114 734 129498 856
rect 129666 734 129958 856
rect 130126 734 130510 856
rect 130678 734 131062 856
rect 131230 734 131522 856
rect 131690 734 132074 856
rect 132242 734 132534 856
rect 132702 734 133086 856
rect 133254 734 133638 856
rect 133806 734 134098 856
rect 134266 734 134650 856
rect 134818 734 135202 856
rect 135370 734 135662 856
rect 135830 734 136214 856
rect 136382 734 136674 856
rect 136842 734 137226 856
rect 137394 734 137778 856
rect 137946 734 138238 856
rect 138406 734 138790 856
rect 138958 734 139250 856
rect 139418 734 139802 856
rect 139970 734 140354 856
rect 140522 734 140814 856
rect 140982 734 141366 856
rect 141534 734 141826 856
rect 141994 734 142378 856
rect 142546 734 142930 856
rect 143098 734 143390 856
rect 143558 734 143942 856
rect 144110 734 144402 856
rect 144570 734 144954 856
rect 145122 734 145506 856
rect 145674 734 145966 856
rect 146134 734 146518 856
rect 146686 734 146978 856
rect 147146 734 147530 856
rect 147698 734 148082 856
rect 148250 734 148542 856
rect 148710 734 149094 856
rect 149262 734 149554 856
rect 149722 734 150106 856
rect 150274 734 150658 856
rect 150826 734 151118 856
rect 151286 734 151670 856
rect 151838 734 152130 856
rect 152298 734 152682 856
rect 152850 734 153234 856
rect 153402 734 153694 856
rect 153862 734 154246 856
rect 154414 734 154706 856
rect 154874 734 155258 856
rect 155426 734 155810 856
rect 155978 734 156270 856
rect 156438 734 156822 856
rect 156990 734 157282 856
rect 157450 734 157834 856
rect 158002 734 158386 856
rect 158554 734 158846 856
rect 159014 734 159398 856
rect 159566 734 159858 856
rect 160026 734 160410 856
rect 160578 734 160962 856
rect 161130 734 161422 856
rect 161590 734 161974 856
rect 162142 734 162434 856
rect 162602 734 162986 856
rect 163154 734 163538 856
rect 163706 734 163998 856
rect 164166 734 164550 856
rect 164718 734 165010 856
rect 165178 734 165562 856
rect 165730 734 166114 856
rect 166282 734 166574 856
rect 166742 734 167126 856
rect 167294 734 167678 856
rect 167846 734 168138 856
rect 168306 734 168690 856
rect 168858 734 169150 856
rect 169318 734 169702 856
rect 169870 734 170254 856
rect 170422 734 170714 856
rect 170882 734 171266 856
rect 171434 734 171726 856
rect 171894 734 172278 856
rect 172446 734 172830 856
rect 172998 734 173290 856
rect 173458 734 173842 856
rect 174010 734 174302 856
rect 174470 734 174854 856
rect 175022 734 175406 856
rect 175574 734 175866 856
rect 176034 734 176418 856
rect 176586 734 176878 856
rect 177046 734 177430 856
rect 177598 734 177982 856
rect 178150 734 178442 856
rect 178610 734 178994 856
rect 179162 734 179454 856
rect 179622 734 180006 856
rect 180174 734 180558 856
rect 180726 734 181018 856
rect 181186 734 181570 856
rect 181738 734 182030 856
rect 182198 734 182582 856
rect 182750 734 183134 856
rect 183302 734 183594 856
rect 183762 734 184146 856
rect 184314 734 184606 856
rect 184774 734 185158 856
rect 185326 734 185710 856
rect 185878 734 186170 856
rect 186338 734 186722 856
rect 186890 734 187182 856
rect 187350 734 187734 856
rect 187902 734 188286 856
rect 188454 734 188746 856
rect 188914 734 189298 856
rect 189466 734 189758 856
rect 189926 734 190310 856
rect 190478 734 190862 856
rect 191030 734 191322 856
rect 191490 734 191874 856
rect 192042 734 192334 856
rect 192502 734 192886 856
rect 193054 734 193438 856
rect 193606 734 193898 856
rect 194066 734 194450 856
rect 194618 734 194910 856
rect 195078 734 195462 856
rect 195630 734 196014 856
rect 196182 734 196474 856
rect 196642 734 197026 856
rect 197194 734 197486 856
rect 197654 734 198038 856
rect 198206 734 198590 856
rect 198758 734 199050 856
rect 199218 734 199602 856
<< metal3 >>
rect 0 174904 800 175024
rect 199200 174904 200000 175024
rect 0 164840 800 164960
rect 199200 164840 200000 164960
rect 0 154912 800 155032
rect 199200 154912 200000 155032
rect 0 144848 800 144968
rect 199200 144848 200000 144968
rect 0 134920 800 135040
rect 199200 134920 200000 135040
rect 0 124856 800 124976
rect 199200 124856 200000 124976
rect 0 114928 800 115048
rect 199200 114928 200000 115048
rect 0 104864 800 104984
rect 199200 104864 200000 104984
rect 0 94936 800 95056
rect 199200 94936 200000 95056
rect 0 84872 800 84992
rect 199200 84872 200000 84992
rect 0 74808 800 74928
rect 199200 74808 200000 74928
rect 0 64880 800 65000
rect 199200 64880 200000 65000
rect 0 54816 800 54936
rect 199200 54816 200000 54936
rect 0 44888 800 45008
rect 199200 44888 200000 45008
rect 0 34824 800 34944
rect 199200 34824 200000 34944
rect 0 24896 800 25016
rect 199200 24896 200000 25016
rect 0 14832 800 14952
rect 199200 14832 200000 14952
rect 0 4904 800 5024
rect 199200 4904 200000 5024
<< obsm3 >>
rect 800 175104 199200 177377
rect 880 174824 199120 175104
rect 800 165040 199200 174824
rect 880 164760 199120 165040
rect 800 155112 199200 164760
rect 880 154832 199120 155112
rect 800 145048 199200 154832
rect 880 144768 199120 145048
rect 800 135120 199200 144768
rect 880 134840 199120 135120
rect 800 125056 199200 134840
rect 880 124776 199120 125056
rect 800 115128 199200 124776
rect 880 114848 199120 115128
rect 800 105064 199200 114848
rect 880 104784 199120 105064
rect 800 95136 199200 104784
rect 880 94856 199120 95136
rect 800 85072 199200 94856
rect 880 84792 199120 85072
rect 800 75008 199200 84792
rect 880 74728 199120 75008
rect 800 65080 199200 74728
rect 880 64800 199120 65080
rect 800 55016 199200 64800
rect 880 54736 199120 55016
rect 800 45088 199200 54736
rect 880 44808 199120 45088
rect 800 35024 199200 44808
rect 880 34744 199120 35024
rect 800 25096 199200 34744
rect 880 24816 199120 25096
rect 800 15032 199200 24816
rect 880 14752 199120 15032
rect 800 5104 199200 14752
rect 880 4824 199120 5104
rect 800 2143 199200 4824
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
rect 188528 2128 188848 177392
<< obsm4 >>
rect 39803 3163 50208 176901
rect 50688 3163 65568 176901
rect 66048 3163 80928 176901
rect 81408 3163 87341 176901
<< labels >>
rlabel metal3 s 199200 4904 200000 5024 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 167826 179200 167882 180000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 160190 179200 160246 180000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 152462 179200 152518 180000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 144734 179200 144790 180000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 137098 179200 137154 180000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 129370 179200 129426 180000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 121642 179200 121698 180000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 114006 179200 114062 180000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 106278 179200 106334 180000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 98642 179200 98698 180000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 199200 34824 200000 34944 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 90914 179200 90970 180000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 83186 179200 83242 180000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 75550 179200 75606 180000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 67822 179200 67878 180000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 60186 179200 60242 180000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 52458 179200 52514 180000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 44730 179200 44786 180000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 37094 179200 37150 180000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 29366 179200 29422 180000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 21638 179200 21694 180000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 199200 64880 200000 65000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 14002 179200 14058 180000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 6274 179200 6330 180000 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 154912 800 155032 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 64880 800 65000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 199200 94936 200000 95056 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 199200 124856 200000 124976 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 199200 154912 200000 155032 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 198646 179200 198702 180000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 190918 179200 190974 180000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 183190 179200 183246 180000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 175554 179200 175610 180000 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 199200 24896 200000 25016 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 162674 179200 162730 180000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 155038 179200 155094 180000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 147310 179200 147366 180000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 139674 179200 139730 180000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 131946 179200 132002 180000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 124218 179200 124274 180000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 116582 179200 116638 180000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 108854 179200 108910 180000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 101218 179200 101274 180000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 93490 179200 93546 180000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 199200 54816 200000 54936 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 85762 179200 85818 180000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 78126 179200 78182 180000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70398 179200 70454 180000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 62670 179200 62726 180000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 55034 179200 55090 180000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 47306 179200 47362 180000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 39670 179200 39726 180000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 31942 179200 31998 180000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 24214 179200 24270 180000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 16578 179200 16634 180000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 199200 84872 200000 84992 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 8850 179200 8906 180000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 1214 179200 1270 180000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 174904 800 175024 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 199200 114928 200000 115048 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 199200 144848 200000 144968 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 199200 174904 200000 175024 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 193494 179200 193550 180000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 185766 179200 185822 180000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 178130 179200 178186 180000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 170402 179200 170458 180000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 199200 14832 200000 14952 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 165250 179200 165306 180000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 157614 179200 157670 180000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 149886 179200 149942 180000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 142158 179200 142214 180000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 134522 179200 134578 180000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 126794 179200 126850 180000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 119158 179200 119214 180000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 111430 179200 111486 180000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 103702 179200 103758 180000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 96066 179200 96122 180000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 199200 44888 200000 45008 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 88338 179200 88394 180000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 80702 179200 80758 180000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 72974 179200 73030 180000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 65246 179200 65302 180000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 57610 179200 57666 180000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 49882 179200 49938 180000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42154 179200 42210 180000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 34518 179200 34574 180000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 26790 179200 26846 180000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 19154 179200 19210 180000 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 199200 74808 200000 74928 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 11426 179200 11482 180000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 3698 179200 3754 180000 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 164840 800 164960 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 104864 800 104984 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 199200 104864 200000 104984 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 199200 134920 200000 135040 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 199200 164840 200000 164960 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 196070 179200 196126 180000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 188342 179200 188398 180000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 180706 179200 180762 180000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 172978 179200 173034 180000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 187238 0 187294 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 102230 0 102286 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 202 0 258 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 170770 0 170826 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 181626 0 181682 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 184662 0 184718 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 186226 0 186282 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 187790 0 187846 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 192390 0 192446 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 193954 0 194010 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 84198 0 84254 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 90362 0 90418 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 91926 0 91982 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 96526 0 96582 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 104254 0 104310 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 153750 0 153806 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 662 0 718 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 183650 0 183706 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 user_clock2
port 502 nsew signal input
rlabel metal4 s 4208 2128 4528 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 34928 2128 35248 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 65648 2128 65968 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 96368 2128 96688 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 127088 2128 127408 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 157808 2128 158128 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 188528 2128 188848 177392 6 vccd1
port 503 nsew power input
rlabel metal4 s 19568 2128 19888 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 50288 2128 50608 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 81008 2128 81328 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 111728 2128 112048 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 142448 2128 142768 177392 6 vssd1
port 504 nsew ground input
rlabel metal4 s 173168 2128 173488 177392 6 vssd1
port 504 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 200000 180000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16527476
string GDS_FILE /home/jasteve4/Documents/ActuatorController/openlane/braille_driver_controller/runs/braille_driver_controller/results/finishing/braille_driver_controller.magic.gds
string GDS_START 799348
<< end >>

