magic
tech sky130A
magscale 1 2
timestamp 1647482984
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 292574 700884 292580 700936
rect 292632 700924 292638 700936
rect 332502 700924 332508 700936
rect 292632 700896 332508 700924
rect 292632 700884 292638 700896
rect 332502 700884 332508 700896
rect 332560 700884 332566 700936
rect 295334 700816 295340 700868
rect 295392 700856 295398 700868
rect 348786 700856 348792 700868
rect 295392 700828 348792 700856
rect 295392 700816 295398 700828
rect 348786 700816 348792 700828
rect 348844 700816 348850 700868
rect 298094 700748 298100 700800
rect 298152 700788 298158 700800
rect 364978 700788 364984 700800
rect 298152 700760 364984 700788
rect 298152 700748 298158 700760
rect 364978 700748 364984 700760
rect 365036 700748 365042 700800
rect 300854 700680 300860 700732
rect 300912 700720 300918 700732
rect 397454 700720 397460 700732
rect 300912 700692 397460 700720
rect 300912 700680 300918 700692
rect 397454 700680 397460 700692
rect 397512 700680 397518 700732
rect 302234 700612 302240 700664
rect 302292 700652 302298 700664
rect 413646 700652 413652 700664
rect 302292 700624 413652 700652
rect 302292 700612 302298 700624
rect 413646 700612 413652 700624
rect 413704 700612 413710 700664
rect 304994 700544 305000 700596
rect 305052 700584 305058 700596
rect 429838 700584 429844 700596
rect 305052 700556 429844 700584
rect 305052 700544 305058 700556
rect 429838 700544 429844 700556
rect 429896 700544 429902 700596
rect 307754 700476 307760 700528
rect 307812 700516 307818 700528
rect 462314 700516 462320 700528
rect 307812 700488 462320 700516
rect 307812 700476 307818 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 310514 700408 310520 700460
rect 310572 700448 310578 700460
rect 478506 700448 478512 700460
rect 310572 700420 478512 700448
rect 310572 700408 310578 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 316034 700340 316040 700392
rect 316092 700380 316098 700392
rect 527174 700380 527180 700392
rect 316092 700352 527180 700380
rect 316092 700340 316098 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 170306 700272 170312 700324
rect 170364 700312 170370 700324
rect 192478 700312 192484 700324
rect 170364 700284 192484 700312
rect 170364 700272 170370 700284
rect 192478 700272 192484 700284
rect 192536 700272 192542 700324
rect 202782 700272 202788 700324
rect 202840 700312 202846 700324
rect 220078 700312 220084 700324
rect 202840 700284 220084 700312
rect 202840 700272 202846 700284
rect 220078 700272 220084 700284
rect 220136 700272 220142 700324
rect 235166 700272 235172 700324
rect 235224 700312 235230 700324
rect 282178 700312 282184 700324
rect 235224 700284 282184 700312
rect 235224 700272 235230 700284
rect 282178 700272 282184 700284
rect 282236 700272 282242 700324
rect 291838 700272 291844 700324
rect 291896 700312 291902 700324
rect 300118 700312 300124 700324
rect 291896 700284 300124 700312
rect 291896 700272 291902 700284
rect 300118 700272 300124 700284
rect 300176 700272 300182 700324
rect 318794 700272 318800 700324
rect 318852 700312 318858 700324
rect 543458 700312 543464 700324
rect 318852 700284 543464 700312
rect 318852 700272 318858 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 283834 700068 283840 700120
rect 283892 700108 283898 700120
rect 284938 700108 284944 700120
rect 283892 700080 284944 700108
rect 283892 700068 283898 700080
rect 284938 700068 284944 700080
rect 284996 700068 285002 700120
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 322934 696940 322940 696992
rect 322992 696980 322998 696992
rect 580166 696980 580172 696992
rect 322992 696952 580172 696980
rect 322992 696940 322998 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 93118 683176 93124 683188
rect 3476 683148 93124 683176
rect 3476 683136 3482 683148
rect 93118 683136 93124 683148
rect 93176 683136 93182 683188
rect 325694 683136 325700 683188
rect 325752 683176 325758 683188
rect 580166 683176 580172 683188
rect 325752 683148 580172 683176
rect 325752 683136 325758 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 328454 670692 328460 670744
rect 328512 670732 328518 670744
rect 580166 670732 580172 670744
rect 328512 670704 580172 670732
rect 328512 670692 328518 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 246298 656928 246304 656940
rect 3568 656900 246304 656928
rect 3568 656888 3574 656900
rect 246298 656888 246304 656900
rect 246356 656888 246362 656940
rect 331214 643084 331220 643136
rect 331272 643124 331278 643136
rect 580166 643124 580172 643136
rect 331272 643096 580172 643124
rect 331272 643084 331278 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 244274 632108 244280 632120
rect 3568 632080 244280 632108
rect 3568 632068 3574 632080
rect 244274 632068 244280 632080
rect 244332 632068 244338 632120
rect 333974 630640 333980 630692
rect 334032 630680 334038 630692
rect 580166 630680 580172 630692
rect 334032 630652 580172 630680
rect 334032 630640 334038 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 336734 616836 336740 616888
rect 336792 616876 336798 616888
rect 580166 616876 580172 616888
rect 336792 616848 580172 616876
rect 336792 616836 336798 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3326 605820 3332 605872
rect 3384 605860 3390 605872
rect 238018 605860 238024 605872
rect 3384 605832 238024 605860
rect 3384 605820 3390 605832
rect 238018 605820 238024 605832
rect 238076 605820 238082 605872
rect 338114 590656 338120 590708
rect 338172 590696 338178 590708
rect 579798 590696 579804 590708
rect 338172 590668 579804 590696
rect 338172 590656 338178 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 235258 579680 235264 579692
rect 3384 579652 235264 579680
rect 3384 579640 3390 579652
rect 235258 579640 235264 579652
rect 235316 579640 235322 579692
rect 340874 576852 340880 576904
rect 340932 576892 340938 576904
rect 580166 576892 580172 576904
rect 340932 576864 580172 576892
rect 340932 576852 340938 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 343634 563048 343640 563100
rect 343692 563088 343698 563100
rect 579798 563088 579804 563100
rect 343692 563060 579804 563088
rect 343692 563048 343698 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 346394 536800 346400 536852
rect 346452 536840 346458 536852
rect 580166 536840 580172 536852
rect 346452 536812 580172 536840
rect 346452 536800 346458 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 228358 527184 228364 527196
rect 3016 527156 228364 527184
rect 3016 527144 3022 527156
rect 228358 527144 228364 527156
rect 228416 527144 228422 527196
rect 349154 524424 349160 524476
rect 349212 524464 349218 524476
rect 580166 524464 580172 524476
rect 349212 524436 580172 524464
rect 349212 524424 349218 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 226334 514808 226340 514820
rect 3384 514780 226340 514808
rect 3384 514768 3390 514780
rect 226334 514768 226340 514780
rect 226392 514768 226398 514820
rect 351914 510620 351920 510672
rect 351972 510660 351978 510672
rect 580166 510660 580172 510672
rect 351972 510632 580172 510660
rect 351972 510620 351978 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 354674 484372 354680 484424
rect 354732 484412 354738 484424
rect 580166 484412 580172 484424
rect 354732 484384 580172 484412
rect 354732 484372 354738 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 220078 476756 220084 476808
rect 220136 476796 220142 476808
rect 277394 476796 277400 476808
rect 220136 476768 277400 476796
rect 220136 476756 220142 476768
rect 277394 476756 277400 476768
rect 277452 476756 277458 476808
rect 2866 474716 2872 474768
rect 2924 474756 2930 474768
rect 220078 474756 220084 474768
rect 2924 474728 220084 474756
rect 2924 474716 2930 474728
rect 220078 474716 220084 474728
rect 220136 474716 220142 474768
rect 356054 470568 356060 470620
rect 356112 470608 356118 470620
rect 579982 470608 579988 470620
rect 356112 470580 579988 470608
rect 356112 470568 356118 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 358814 456764 358820 456816
rect 358872 456804 358878 456816
rect 580166 456804 580172 456816
rect 358872 456776 580172 456804
rect 358872 456764 358878 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 361574 430584 361580 430636
rect 361632 430624 361638 430636
rect 580166 430624 580172 430636
rect 361632 430596 580172 430624
rect 361632 430584 361638 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 2774 423512 2780 423564
rect 2832 423552 2838 423564
rect 4798 423552 4804 423564
rect 2832 423524 4804 423552
rect 2832 423512 2838 423524
rect 4798 423512 4804 423524
rect 4856 423512 4862 423564
rect 364334 418140 364340 418192
rect 364392 418180 364398 418192
rect 580166 418180 580172 418192
rect 364392 418152 580172 418180
rect 364392 418140 364398 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 3326 409844 3332 409896
rect 3384 409884 3390 409896
rect 211154 409884 211160 409896
rect 3384 409856 211160 409884
rect 3384 409844 3390 409856
rect 211154 409844 211160 409856
rect 211212 409844 211218 409896
rect 367094 404336 367100 404388
rect 367152 404376 367158 404388
rect 580166 404376 580172 404388
rect 367152 404348 580172 404376
rect 367152 404336 367158 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 369854 378156 369860 378208
rect 369912 378196 369918 378208
rect 580166 378196 580172 378208
rect 369912 378168 580172 378196
rect 369912 378156 369918 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 136634 371832 136640 371884
rect 136692 371872 136698 371884
rect 269666 371872 269672 371884
rect 136692 371844 269672 371872
rect 136692 371832 136698 371844
rect 269666 371832 269672 371844
rect 269724 371832 269730 371884
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 13814 371260 13820 371272
rect 3384 371232 13820 371260
rect 3384 371220 3390 371232
rect 13814 371220 13820 371232
rect 13872 371220 13878 371272
rect 93118 370472 93124 370524
rect 93176 370512 93182 370524
rect 251818 370512 251824 370524
rect 93176 370484 251824 370512
rect 93176 370472 93182 370484
rect 251818 370472 251824 370484
rect 251876 370472 251882 370524
rect 13814 369112 13820 369164
rect 13872 369152 13878 369164
rect 205634 369152 205640 369164
rect 13872 369124 205640 369152
rect 13872 369112 13878 369124
rect 205634 369112 205640 369124
rect 205692 369112 205698 369164
rect 4798 367752 4804 367804
rect 4856 367792 4862 367804
rect 213178 367792 213184 367804
rect 4856 367764 213184 367792
rect 4856 367752 4862 367764
rect 213178 367752 213184 367764
rect 213236 367752 213242 367804
rect 40034 366324 40040 366376
rect 40092 366364 40098 366376
rect 259822 366364 259828 366376
rect 40092 366336 259828 366364
rect 40092 366324 40098 366336
rect 259822 366324 259828 366336
rect 259880 366324 259886 366376
rect 104894 364964 104900 365016
rect 104952 365004 104958 365016
rect 267550 365004 267556 365016
rect 104952 364976 267556 365004
rect 104952 364964 104958 364976
rect 267550 364964 267556 364976
rect 267608 364964 267614 365016
rect 372706 364352 372712 364404
rect 372764 364392 372770 364404
rect 580166 364392 580172 364404
rect 372764 364364 580172 364392
rect 372764 364352 372770 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 192478 363604 192484 363656
rect 192536 363644 192542 363656
rect 275186 363644 275192 363656
rect 192536 363616 275192 363644
rect 192536 363604 192542 363616
rect 275186 363604 275192 363616
rect 275244 363604 275250 363656
rect 228358 363196 228364 363248
rect 228416 363236 228422 363248
rect 229094 363236 229100 363248
rect 228416 363208 229100 363236
rect 228416 363196 228422 363208
rect 229094 363196 229100 363208
rect 229152 363196 229158 363248
rect 238018 363196 238024 363248
rect 238076 363236 238082 363248
rect 239306 363236 239312 363248
rect 238076 363208 239312 363236
rect 238076 363196 238082 363208
rect 239306 363196 239312 363208
rect 239364 363196 239370 363248
rect 220078 362924 220084 362976
rect 220136 362964 220142 362976
rect 221366 362964 221372 362976
rect 220136 362936 221372 362964
rect 220136 362924 220142 362936
rect 221366 362924 221372 362936
rect 221424 362924 221430 362976
rect 235258 362924 235264 362976
rect 235316 362964 235322 362976
rect 236730 362964 236736 362976
rect 235316 362936 236736 362964
rect 235316 362924 235322 362936
rect 236730 362924 236736 362936
rect 236788 362924 236794 362976
rect 246298 362924 246304 362976
rect 246356 362964 246362 362976
rect 247034 362964 247040 362976
rect 246356 362936 247040 362964
rect 246356 362924 246362 362936
rect 247034 362924 247040 362936
rect 247092 362924 247098 362976
rect 71774 362856 71780 362908
rect 71832 362896 71838 362908
rect 262398 362896 262404 362908
rect 71832 362868 262404 362896
rect 71832 362856 71838 362868
rect 262398 362856 262404 362868
rect 262456 362856 262462 362908
rect 284938 362856 284944 362908
rect 284996 362896 285002 362908
rect 288066 362896 288072 362908
rect 284996 362868 288072 362896
rect 284996 362856 285002 362868
rect 288066 362856 288072 362868
rect 288124 362856 288130 362908
rect 4062 362788 4068 362840
rect 4120 362828 4126 362840
rect 208578 362828 208584 362840
rect 4120 362800 208584 362828
rect 4120 362788 4126 362800
rect 208578 362788 208584 362800
rect 208636 362788 208642 362840
rect 218054 362788 218060 362840
rect 218112 362828 218118 362840
rect 280338 362828 280344 362840
rect 218112 362800 280344 362828
rect 218112 362788 218118 362800
rect 280338 362788 280344 362800
rect 280396 362788 280402 362840
rect 3970 362720 3976 362772
rect 4028 362760 4034 362772
rect 216214 362760 216220 362772
rect 4028 362732 216220 362760
rect 4028 362720 4034 362732
rect 216214 362720 216220 362732
rect 216272 362720 216278 362772
rect 3878 362652 3884 362704
rect 3936 362692 3942 362704
rect 218790 362692 218796 362704
rect 3936 362664 218796 362692
rect 3936 362652 3942 362664
rect 218790 362652 218796 362664
rect 218848 362652 218854 362704
rect 3786 362584 3792 362636
rect 3844 362624 3850 362636
rect 223942 362624 223948 362636
rect 3844 362596 223948 362624
rect 3844 362584 3850 362596
rect 223942 362584 223948 362596
rect 224000 362584 224006 362636
rect 3694 362516 3700 362568
rect 3752 362556 3758 362568
rect 231670 362556 231676 362568
rect 3752 362528 231676 362556
rect 3752 362516 3758 362528
rect 231670 362516 231676 362528
rect 231728 362516 231734 362568
rect 3602 362448 3608 362500
rect 3660 362488 3666 362500
rect 234154 362488 234160 362500
rect 3660 362460 234160 362488
rect 3660 362448 3666 362460
rect 234154 362448 234160 362460
rect 234212 362448 234218 362500
rect 23474 362380 23480 362432
rect 23532 362420 23538 362432
rect 257246 362420 257252 362432
rect 23532 362392 257252 362420
rect 23532 362380 23538 362392
rect 257246 362380 257252 362392
rect 257304 362380 257310 362432
rect 3510 362312 3516 362364
rect 3568 362352 3574 362364
rect 241882 362352 241888 362364
rect 3568 362324 241888 362352
rect 3568 362312 3574 362324
rect 241882 362312 241888 362324
rect 241940 362312 241946 362364
rect 3418 362244 3424 362296
rect 3476 362284 3482 362296
rect 249610 362284 249616 362296
rect 3476 362256 249616 362284
rect 3476 362244 3482 362256
rect 249610 362244 249616 362256
rect 249668 362244 249674 362296
rect 313642 362244 313648 362296
rect 313700 362284 313706 362296
rect 494054 362284 494060 362296
rect 313700 362256 494060 362284
rect 313700 362244 313706 362256
rect 494054 362244 494060 362256
rect 494112 362244 494118 362296
rect 6914 362176 6920 362228
rect 6972 362216 6978 362228
rect 254670 362216 254676 362228
rect 6972 362188 254676 362216
rect 6972 362176 6978 362188
rect 254670 362176 254676 362188
rect 254728 362176 254734 362228
rect 266354 362176 266360 362228
rect 266412 362216 266418 362228
rect 285490 362216 285496 362228
rect 266412 362188 285496 362216
rect 266412 362176 266418 362188
rect 285490 362176 285496 362188
rect 285548 362176 285554 362228
rect 321370 362176 321376 362228
rect 321428 362216 321434 362228
rect 558914 362216 558920 362228
rect 321428 362188 558920 362216
rect 321428 362176 321434 362188
rect 558914 362176 558920 362188
rect 558972 362176 558978 362228
rect 88334 362108 88340 362160
rect 88392 362148 88398 362160
rect 264974 362148 264980 362160
rect 88392 362120 264980 362148
rect 88392 362108 88398 362120
rect 264974 362108 264980 362120
rect 265032 362108 265038 362160
rect 153194 362040 153200 362092
rect 153252 362080 153258 362092
rect 272702 362080 272708 362092
rect 153252 362052 272708 362080
rect 153252 362040 153258 362052
rect 272702 362040 272708 362052
rect 272760 362040 272766 362092
rect 382918 361904 382924 361956
rect 382976 361944 382982 361956
rect 479518 361944 479524 361956
rect 382976 361916 479524 361944
rect 382976 361904 382982 361916
rect 479518 361904 479524 361916
rect 479576 361904 479582 361956
rect 282178 361836 282184 361888
rect 282236 361876 282242 361888
rect 282914 361876 282920 361888
rect 282236 361848 282920 361876
rect 282236 361836 282242 361848
rect 282914 361836 282920 361848
rect 282972 361836 282978 361888
rect 290642 361836 290648 361888
rect 290700 361876 290706 361888
rect 291838 361876 291844 361888
rect 290700 361848 291844 361876
rect 290700 361836 290706 361848
rect 291838 361836 291844 361848
rect 291896 361836 291902 361888
rect 388070 361836 388076 361888
rect 388128 361876 388134 361888
rect 486418 361876 486424 361888
rect 388128 361848 486424 361876
rect 388128 361836 388134 361848
rect 486418 361836 486424 361848
rect 486476 361836 486482 361888
rect 385494 361768 385500 361820
rect 385552 361808 385558 361820
rect 483658 361808 483664 361820
rect 385552 361780 483664 361808
rect 385552 361768 385558 361780
rect 483658 361768 483664 361780
rect 483716 361768 483722 361820
rect 377766 361700 377772 361752
rect 377824 361740 377830 361752
rect 485038 361740 485044 361752
rect 377824 361712 485044 361740
rect 377824 361700 377830 361712
rect 485038 361700 485044 361712
rect 485096 361700 485102 361752
rect 375190 361632 375196 361684
rect 375248 361672 375254 361684
rect 482278 361672 482284 361684
rect 375248 361644 482284 361672
rect 375248 361632 375254 361644
rect 482278 361632 482284 361644
rect 482336 361632 482342 361684
rect 380342 361564 380348 361616
rect 380400 361604 380406 361616
rect 489178 361604 489184 361616
rect 380400 361576 489184 361604
rect 380400 361564 380406 361576
rect 489178 361564 489184 361576
rect 489236 361564 489242 361616
rect 186958 360476 186964 360528
rect 187016 360516 187022 360528
rect 195698 360516 195704 360528
rect 187016 360488 195704 360516
rect 187016 360476 187022 360488
rect 195698 360476 195704 360488
rect 195756 360476 195762 360528
rect 4798 360408 4804 360460
rect 4856 360448 4862 360460
rect 198274 360448 198280 360460
rect 4856 360420 198280 360448
rect 4856 360408 4862 360420
rect 198274 360408 198280 360420
rect 198332 360408 198338 360460
rect 191098 360340 191104 360392
rect 191156 360380 191162 360392
rect 200850 360380 200856 360392
rect 191156 360352 200856 360380
rect 191156 360340 191162 360352
rect 200850 360340 200856 360352
rect 200908 360340 200914 360392
rect 191742 360272 191748 360324
rect 191800 360312 191806 360324
rect 203426 360312 203432 360324
rect 191800 360284 203432 360312
rect 191800 360272 191806 360284
rect 203426 360272 203432 360284
rect 203484 360272 203490 360324
rect 188338 360204 188344 360256
rect 188396 360244 188402 360256
rect 193214 360244 193220 360256
rect 188396 360216 193220 360244
rect 188396 360204 188402 360216
rect 193214 360204 193220 360216
rect 193272 360204 193278 360256
rect 390922 359388 390928 359440
rect 390980 359428 390986 359440
rect 391842 359428 391848 359440
rect 390980 359400 391848 359428
rect 390980 359388 390986 359400
rect 391842 359388 391848 359400
rect 391900 359388 391906 359440
rect 391842 358776 391848 358828
rect 391900 358816 391906 358828
rect 406378 358816 406384 358828
rect 391900 358788 406384 358816
rect 391900 358776 391906 358788
rect 406378 358776 406384 358788
rect 406436 358776 406442 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 191742 358748 191748 358760
rect 3384 358720 191748 358748
rect 3384 358708 3390 358720
rect 191742 358708 191748 358720
rect 191800 358708 191806 358760
rect 482278 353200 482284 353252
rect 482336 353240 482342 353252
rect 580166 353240 580172 353252
rect 482336 353212 580172 353240
rect 482336 353200 482342 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 191098 346372 191104 346384
rect 3200 346344 191104 346372
rect 3200 346332 3206 346344
rect 191098 346332 191104 346344
rect 191156 346332 191162 346384
rect 3418 343612 3424 343664
rect 3476 343652 3482 343664
rect 189074 343652 189080 343664
rect 3476 343624 189080 343652
rect 3476 343612 3482 343624
rect 189074 343612 189080 343624
rect 189132 343612 189138 343664
rect 7558 333956 7564 334008
rect 7616 333996 7622 334008
rect 189074 333996 189080 334008
rect 7616 333968 189080 333996
rect 7616 333956 7622 333968
rect 189074 333956 189080 333968
rect 189132 333956 189138 334008
rect 485038 325592 485044 325644
rect 485096 325632 485102 325644
rect 580166 325632 580172 325644
rect 485096 325604 580172 325632
rect 485096 325592 485102 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 22738 324300 22744 324352
rect 22796 324340 22802 324352
rect 189074 324340 189080 324352
rect 22796 324312 189080 324340
rect 22796 324300 22802 324312
rect 189074 324300 189080 324312
rect 189132 324300 189138 324352
rect 2774 319812 2780 319864
rect 2832 319852 2838 319864
rect 4798 319852 4804 319864
rect 2832 319824 4804 319852
rect 2832 319812 2838 319824
rect 4798 319812 4804 319824
rect 4856 319812 4862 319864
rect 394326 314712 394332 314764
rect 394384 314752 394390 314764
rect 395338 314752 395344 314764
rect 394384 314724 395344 314752
rect 394384 314712 394390 314724
rect 395338 314712 395344 314724
rect 395396 314712 395402 314764
rect 489178 313216 489184 313268
rect 489236 313256 489242 313268
rect 580166 313256 580172 313268
rect 489236 313228 580172 313256
rect 489236 313216 489242 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 186958 306320 186964 306332
rect 3568 306292 186964 306320
rect 3568 306280 3574 306292
rect 186958 306280 186964 306292
rect 187016 306280 187022 306332
rect 4798 303628 4804 303680
rect 4856 303668 4862 303680
rect 189074 303668 189080 303680
rect 4856 303640 189080 303668
rect 4856 303628 4862 303640
rect 189074 303628 189080 303640
rect 189132 303628 189138 303680
rect 394326 303628 394332 303680
rect 394384 303668 394390 303680
rect 554038 303668 554044 303680
rect 394384 303640 554044 303668
rect 394384 303628 394390 303640
rect 554038 303628 554044 303640
rect 554096 303628 554102 303680
rect 479518 299412 479524 299464
rect 479576 299452 479582 299464
rect 580166 299452 580172 299464
rect 479576 299424 580172 299452
rect 479576 299412 479582 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 188338 293944 188344 293956
rect 3108 293916 188344 293944
rect 3108 293904 3114 293916
rect 188338 293904 188344 293916
rect 188396 293904 188402 293956
rect 394418 284520 394424 284572
rect 394476 284560 394482 284572
rect 399478 284560 399484 284572
rect 394476 284532 399484 284560
rect 394476 284520 394482 284532
rect 399478 284520 399484 284532
rect 399536 284520 399542 284572
rect 14458 274660 14464 274712
rect 14516 274700 14522 274712
rect 189074 274700 189080 274712
rect 14516 274672 189080 274700
rect 14516 274660 14522 274672
rect 189074 274660 189080 274672
rect 189132 274660 189138 274712
rect 394418 274660 394424 274712
rect 394476 274700 394482 274712
rect 551278 274700 551284 274712
rect 394476 274672 551284 274700
rect 394476 274660 394482 274672
rect 551278 274660 551284 274672
rect 551336 274660 551342 274712
rect 483658 273164 483664 273216
rect 483716 273204 483722 273216
rect 580166 273204 580172 273216
rect 483716 273176 580172 273204
rect 483716 273164 483722 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3510 267656 3516 267708
rect 3568 267696 3574 267708
rect 7558 267696 7564 267708
rect 3568 267668 7564 267696
rect 3568 267656 3574 267668
rect 7558 267656 7564 267668
rect 7616 267656 7622 267708
rect 486418 259360 486424 259412
rect 486476 259400 486482 259412
rect 580166 259400 580172 259412
rect 486476 259372 580172 259400
rect 486476 259360 486482 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 3602 253920 3608 253972
rect 3660 253960 3666 253972
rect 189074 253960 189080 253972
rect 3660 253932 189080 253960
rect 3660 253920 3666 253932
rect 189074 253920 189080 253932
rect 189132 253920 189138 253972
rect 406378 245556 406384 245608
rect 406436 245596 406442 245608
rect 580166 245596 580172 245608
rect 406436 245568 580172 245596
rect 406436 245556 406442 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 393774 244536 393780 244588
rect 393832 244576 393838 244588
rect 396718 244576 396724 244588
rect 393832 244548 396724 244576
rect 393832 244536 393838 244548
rect 396718 244536 396724 244548
rect 396776 244536 396782 244588
rect 7558 244264 7564 244316
rect 7616 244304 7622 244316
rect 189074 244304 189080 244316
rect 7616 244276 189080 244304
rect 7616 244264 7622 244276
rect 189074 244264 189080 244276
rect 189132 244264 189138 244316
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 189718 241448 189724 241460
rect 3476 241420 189724 241448
rect 3476 241408 3482 241420
rect 189718 241408 189724 241420
rect 189776 241408 189782 241460
rect 394142 233180 394148 233232
rect 394200 233220 394206 233232
rect 579982 233220 579988 233232
rect 394200 233192 579988 233220
rect 394200 233180 394206 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 3510 224952 3516 225004
rect 3568 224992 3574 225004
rect 189074 224992 189080 225004
rect 3568 224964 189080 224992
rect 3568 224952 3574 224964
rect 189074 224952 189080 224964
rect 189132 224952 189138 225004
rect 394050 219376 394056 219428
rect 394108 219416 394114 219428
rect 580166 219416 580172 219428
rect 394108 219388 580172 219416
rect 394108 219376 394114 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 21358 213936 21364 213988
rect 21416 213976 21422 213988
rect 189074 213976 189080 213988
rect 21416 213948 189080 213976
rect 21416 213936 21422 213948
rect 189074 213936 189080 213948
rect 189132 213936 189138 213988
rect 394050 213936 394056 213988
rect 394108 213976 394114 213988
rect 457438 213976 457444 213988
rect 394108 213948 457444 213976
rect 394108 213936 394114 213948
rect 457438 213936 457444 213948
rect 457496 213936 457502 213988
rect 393958 206932 393964 206984
rect 394016 206972 394022 206984
rect 579798 206972 579804 206984
rect 394016 206944 579804 206972
rect 394016 206932 394022 206944
rect 579798 206932 579804 206944
rect 579856 206932 579862 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 190086 202824 190092 202836
rect 3108 202796 190092 202824
rect 3108 202784 3114 202796
rect 190086 202784 190092 202796
rect 190144 202784 190150 202836
rect 3418 194556 3424 194608
rect 3476 194596 3482 194608
rect 189074 194596 189080 194608
rect 3476 194568 189080 194596
rect 3476 194556 3482 194568
rect 189074 194556 189080 194568
rect 189132 194556 189138 194608
rect 394602 193128 394608 193180
rect 394660 193168 394666 193180
rect 580166 193168 580172 193180
rect 394660 193140 580172 193168
rect 394660 193128 394666 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 22738 189020 22744 189032
rect 3200 188992 22744 189020
rect 3200 188980 3206 188992
rect 22738 188980 22744 188992
rect 22796 188980 22802 189032
rect 394602 184900 394608 184952
rect 394660 184940 394666 184952
rect 576118 184940 576124 184952
rect 394660 184912 576124 184940
rect 394660 184900 394666 184912
rect 576118 184900 576124 184912
rect 576176 184900 576182 184952
rect 395338 179324 395344 179376
rect 395396 179364 395402 179376
rect 580166 179364 580172 179376
rect 395396 179336 580172 179364
rect 395396 179324 395402 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 308214 177760 308220 177812
rect 308272 177800 308278 177812
rect 338758 177800 338764 177812
rect 308272 177772 338764 177800
rect 308272 177760 308278 177772
rect 338758 177760 338764 177772
rect 338816 177760 338822 177812
rect 320082 177692 320088 177744
rect 320140 177732 320146 177744
rect 418154 177732 418160 177744
rect 320140 177704 418160 177732
rect 320140 177692 320146 177704
rect 418154 177692 418160 177704
rect 418212 177692 418218 177744
rect 188338 177624 188344 177676
rect 188396 177664 188402 177676
rect 203702 177664 203708 177676
rect 188396 177636 203708 177664
rect 188396 177624 188402 177636
rect 203702 177624 203708 177636
rect 203760 177624 203766 177676
rect 209314 177624 209320 177676
rect 209372 177664 209378 177676
rect 224954 177664 224960 177676
rect 209372 177636 224960 177664
rect 209372 177624 209378 177636
rect 224954 177624 224960 177636
rect 225012 177624 225018 177676
rect 323210 177624 323216 177676
rect 323268 177664 323274 177676
rect 425054 177664 425060 177676
rect 323268 177636 425060 177664
rect 323268 177624 323274 177636
rect 425054 177624 425060 177636
rect 425112 177624 425118 177676
rect 191098 177556 191104 177608
rect 191156 177596 191162 177608
rect 211430 177596 211436 177608
rect 191156 177568 211436 177596
rect 191156 177556 191162 177568
rect 211430 177556 211436 177568
rect 211488 177556 211494 177608
rect 227898 177556 227904 177608
rect 227956 177596 227962 177608
rect 236638 177596 236644 177608
rect 227956 177568 236644 177596
rect 227956 177556 227962 177568
rect 236638 177556 236644 177568
rect 236696 177556 236702 177608
rect 326522 177556 326528 177608
rect 326580 177596 326586 177608
rect 431954 177596 431960 177608
rect 326580 177568 431960 177596
rect 326580 177556 326586 177568
rect 431954 177556 431960 177568
rect 432012 177556 432018 177608
rect 184934 177488 184940 177540
rect 184992 177528 184998 177540
rect 217134 177528 217140 177540
rect 184992 177500 217140 177528
rect 184992 177488 184998 177500
rect 217134 177488 217140 177500
rect 217192 177488 217198 177540
rect 248230 177488 248236 177540
rect 248288 177528 248294 177540
rect 251818 177528 251824 177540
rect 248288 177500 251824 177528
rect 248288 177488 248294 177500
rect 251818 177488 251824 177500
rect 251876 177488 251882 177540
rect 262214 177488 262220 177540
rect 262272 177488 262278 177540
rect 265250 177488 265256 177540
rect 265308 177528 265314 177540
rect 282178 177528 282184 177540
rect 265308 177500 282184 177528
rect 265308 177488 265314 177500
rect 282178 177488 282184 177500
rect 282236 177488 282242 177540
rect 290182 177488 290188 177540
rect 290240 177528 290246 177540
rect 300026 177528 300032 177540
rect 290240 177500 300032 177528
rect 290240 177488 290246 177500
rect 300026 177488 300032 177500
rect 300084 177488 300090 177540
rect 300854 177488 300860 177540
rect 300912 177528 300918 177540
rect 309962 177528 309968 177540
rect 300912 177500 309968 177528
rect 300912 177488 300918 177500
rect 309962 177488 309968 177500
rect 310020 177488 310026 177540
rect 329650 177488 329656 177540
rect 329708 177528 329714 177540
rect 440234 177528 440240 177540
rect 329708 177500 440240 177528
rect 329708 177488 329714 177500
rect 440234 177488 440240 177500
rect 440292 177488 440298 177540
rect 176654 177420 176660 177472
rect 176712 177460 176718 177472
rect 214006 177460 214012 177472
rect 176712 177432 214012 177460
rect 176712 177420 176718 177432
rect 214006 177420 214012 177432
rect 214064 177420 214070 177472
rect 214558 177420 214564 177472
rect 214616 177460 214622 177472
rect 225782 177460 225788 177472
rect 214616 177432 225788 177460
rect 214616 177420 214622 177432
rect 225782 177420 225788 177432
rect 225840 177420 225846 177472
rect 248138 177420 248144 177472
rect 248196 177460 248202 177472
rect 252554 177460 252560 177472
rect 248196 177432 252560 177460
rect 248196 177420 248202 177432
rect 252554 177420 252560 177432
rect 252612 177420 252618 177472
rect 262232 177460 262260 177488
rect 285674 177460 285680 177472
rect 262232 177432 285680 177460
rect 285674 177420 285680 177432
rect 285732 177420 285738 177472
rect 286226 177420 286232 177472
rect 286284 177460 286290 177472
rect 307018 177460 307024 177472
rect 286284 177432 307024 177460
rect 286284 177420 286290 177432
rect 307018 177420 307024 177432
rect 307076 177420 307082 177472
rect 332502 177420 332508 177472
rect 332560 177460 332566 177472
rect 447134 177460 447140 177472
rect 332560 177432 447140 177460
rect 332560 177420 332566 177432
rect 447134 177420 447140 177432
rect 447192 177420 447198 177472
rect 141418 177352 141424 177404
rect 141476 177392 141482 177404
rect 195422 177392 195428 177404
rect 141476 177364 195428 177392
rect 141476 177352 141482 177364
rect 195422 177352 195428 177364
rect 195480 177352 195486 177404
rect 206278 177352 206284 177404
rect 206336 177392 206342 177404
rect 226886 177392 226892 177404
rect 206336 177364 226892 177392
rect 206336 177352 206342 177364
rect 226886 177352 226892 177364
rect 226944 177352 226950 177404
rect 246206 177352 246212 177404
rect 246264 177392 246270 177404
rect 250070 177392 250076 177404
rect 246264 177364 250076 177392
rect 246264 177352 246270 177364
rect 250070 177352 250076 177364
rect 250128 177352 250134 177404
rect 252186 177352 252192 177404
rect 252244 177392 252250 177404
rect 262214 177392 262220 177404
rect 252244 177364 262220 177392
rect 252244 177352 252250 177364
rect 262214 177352 262220 177364
rect 262272 177352 262278 177404
rect 264514 177352 264520 177404
rect 264572 177392 264578 177404
rect 291194 177392 291200 177404
rect 264572 177364 291200 177392
rect 264572 177352 264578 177364
rect 291194 177352 291200 177364
rect 291252 177352 291258 177404
rect 302142 177352 302148 177404
rect 302200 177392 302206 177404
rect 312538 177392 312544 177404
rect 302200 177364 312544 177392
rect 302200 177352 302206 177364
rect 312538 177352 312544 177364
rect 312596 177352 312602 177404
rect 315942 177352 315948 177404
rect 316000 177392 316006 177404
rect 320818 177392 320824 177404
rect 316000 177364 320824 177392
rect 316000 177352 316006 177364
rect 320818 177352 320824 177364
rect 320876 177352 320882 177404
rect 335354 177352 335360 177404
rect 335412 177392 335418 177404
rect 454034 177392 454040 177404
rect 335412 177364 454040 177392
rect 335412 177352 335418 177364
rect 454034 177352 454040 177364
rect 454092 177352 454098 177404
rect 134518 177284 134524 177336
rect 134576 177324 134582 177336
rect 192294 177324 192300 177336
rect 134576 177296 192300 177324
rect 134576 177284 134582 177296
rect 192294 177284 192300 177296
rect 192352 177284 192358 177336
rect 201494 177284 201500 177336
rect 201552 177324 201558 177336
rect 225414 177324 225420 177336
rect 201552 177296 225420 177324
rect 201552 177284 201558 177296
rect 225414 177284 225420 177296
rect 225472 177284 225478 177336
rect 247586 177284 247592 177336
rect 247644 177324 247650 177336
rect 251266 177324 251272 177336
rect 247644 177296 251272 177324
rect 247644 177284 247650 177296
rect 251266 177284 251272 177296
rect 251324 177284 251330 177336
rect 252370 177284 252376 177336
rect 252428 177324 252434 177336
rect 263594 177324 263600 177336
rect 252428 177296 263600 177324
rect 252428 177284 252434 177296
rect 263594 177284 263600 177296
rect 263652 177284 263658 177336
rect 281718 177284 281724 177336
rect 281776 177324 281782 177336
rect 329098 177324 329104 177336
rect 281776 177296 329104 177324
rect 281776 177284 281782 177296
rect 329098 177284 329104 177296
rect 329156 177284 329162 177336
rect 338482 177284 338488 177336
rect 338540 177324 338546 177336
rect 460934 177324 460940 177336
rect 338540 177296 460940 177324
rect 338540 177284 338546 177296
rect 460934 177284 460940 177296
rect 460992 177284 460998 177336
rect 246114 177216 246120 177268
rect 246172 177256 246178 177268
rect 248414 177256 248420 177268
rect 246172 177228 248420 177256
rect 246172 177216 246178 177228
rect 248414 177216 248420 177228
rect 248472 177216 248478 177268
rect 343634 177148 343640 177200
rect 343692 177188 343698 177200
rect 346946 177188 346952 177200
rect 343692 177160 346952 177188
rect 343692 177148 343698 177160
rect 346946 177148 346952 177160
rect 347004 177148 347010 177200
rect 333146 177080 333152 177132
rect 333204 177120 333210 177132
rect 336182 177120 336188 177132
rect 333204 177092 336188 177120
rect 333204 177080 333210 177092
rect 336182 177080 336188 177092
rect 336240 177080 336246 177132
rect 373718 177012 373724 177064
rect 373776 177052 373782 177064
rect 374638 177052 374644 177064
rect 373776 177024 374644 177052
rect 373776 177012 373782 177024
rect 374638 177012 374644 177024
rect 374696 177012 374702 177064
rect 226334 176944 226340 176996
rect 226392 176984 226398 176996
rect 229186 176984 229192 176996
rect 226392 176956 229192 176984
rect 226392 176944 226398 176956
rect 229186 176944 229192 176956
rect 229244 176944 229250 176996
rect 238018 176944 238024 176996
rect 238076 176984 238082 176996
rect 238846 176984 238852 176996
rect 238076 176956 238852 176984
rect 238076 176944 238082 176956
rect 238846 176944 238852 176956
rect 238904 176944 238910 176996
rect 284202 176944 284208 176996
rect 284260 176984 284266 176996
rect 287698 176984 287704 176996
rect 284260 176956 287704 176984
rect 284260 176944 284266 176956
rect 287698 176944 287704 176956
rect 287756 176944 287762 176996
rect 217594 176876 217600 176928
rect 217652 176916 217658 176928
rect 221182 176916 221188 176928
rect 217652 176888 221188 176916
rect 217652 176876 217658 176888
rect 221182 176876 221188 176888
rect 221240 176876 221246 176928
rect 234706 176876 234712 176928
rect 234764 176916 234770 176928
rect 240226 176916 240232 176928
rect 234764 176888 240232 176916
rect 234764 176876 234770 176888
rect 240226 176876 240232 176888
rect 240284 176876 240290 176928
rect 262122 176876 262128 176928
rect 262180 176916 262186 176928
rect 269666 176916 269672 176928
rect 262180 176888 269672 176916
rect 262180 176876 262186 176888
rect 269666 176876 269672 176888
rect 269724 176876 269730 176928
rect 273162 176876 273168 176928
rect 273220 176916 273226 176928
rect 278038 176916 278044 176928
rect 273220 176888 278044 176916
rect 273220 176876 273226 176888
rect 278038 176876 278044 176888
rect 278096 176876 278102 176928
rect 236270 176808 236276 176860
rect 236328 176848 236334 176860
rect 240318 176848 240324 176860
rect 236328 176820 240324 176848
rect 236328 176808 236334 176820
rect 240318 176808 240324 176820
rect 240376 176808 240382 176860
rect 192478 176672 192484 176724
rect 192536 176712 192542 176724
rect 193398 176712 193404 176724
rect 192536 176684 193404 176712
rect 192536 176672 192542 176684
rect 193398 176672 193404 176684
rect 193456 176672 193462 176724
rect 226978 176672 226984 176724
rect 227036 176712 227042 176724
rect 227806 176712 227812 176724
rect 227036 176684 227812 176712
rect 227036 176672 227042 176684
rect 227806 176672 227812 176684
rect 227864 176672 227870 176724
rect 235258 176672 235264 176724
rect 235316 176712 235322 176724
rect 238294 176712 238300 176724
rect 235316 176684 238300 176712
rect 235316 176672 235322 176684
rect 238294 176672 238300 176684
rect 238352 176672 238358 176724
rect 240778 176672 240784 176724
rect 240836 176712 240842 176724
rect 241514 176712 241520 176724
rect 240836 176684 241520 176712
rect 240836 176672 240842 176684
rect 241514 176672 241520 176684
rect 241572 176672 241578 176724
rect 244826 176672 244832 176724
rect 244884 176712 244890 176724
rect 245746 176712 245752 176724
rect 244884 176684 245752 176712
rect 244884 176672 244890 176684
rect 245746 176672 245752 176684
rect 245804 176672 245810 176724
rect 272978 176672 272984 176724
rect 273036 176712 273042 176724
rect 273898 176712 273904 176724
rect 273036 176684 273904 176712
rect 273036 176672 273042 176684
rect 273898 176672 273904 176684
rect 273956 176672 273962 176724
rect 279050 176672 279056 176724
rect 279108 176712 279114 176724
rect 282270 176712 282276 176724
rect 279108 176684 282276 176712
rect 279108 176672 279114 176684
rect 282270 176672 282276 176684
rect 282328 176672 282334 176724
rect 291010 176672 291016 176724
rect 291068 176712 291074 176724
rect 295978 176712 295984 176724
rect 291068 176684 295984 176712
rect 291068 176672 291074 176684
rect 295978 176672 295984 176684
rect 296036 176672 296042 176724
rect 297450 176672 297456 176724
rect 297508 176712 297514 176724
rect 304258 176712 304264 176724
rect 297508 176684 304264 176712
rect 297508 176672 297514 176684
rect 304258 176672 304264 176684
rect 304316 176672 304322 176724
rect 307570 176672 307576 176724
rect 307628 176712 307634 176724
rect 309870 176712 309876 176724
rect 307628 176684 309876 176712
rect 307628 176672 307634 176684
rect 309870 176672 309876 176684
rect 309928 176672 309934 176724
rect 318886 176672 318892 176724
rect 318944 176712 318950 176724
rect 323578 176712 323584 176724
rect 318944 176684 323584 176712
rect 318944 176672 318950 176684
rect 323578 176672 323584 176684
rect 323636 176672 323642 176724
rect 326982 176672 326988 176724
rect 327040 176712 327046 176724
rect 329190 176712 329196 176724
rect 327040 176684 329196 176712
rect 327040 176672 327046 176684
rect 329190 176672 329196 176684
rect 329248 176672 329254 176724
rect 337470 176672 337476 176724
rect 337528 176712 337534 176724
rect 338850 176712 338856 176724
rect 337528 176684 338856 176712
rect 337528 176672 337534 176684
rect 338850 176672 338856 176684
rect 338908 176672 338914 176724
rect 354950 176672 354956 176724
rect 355008 176712 355014 176724
rect 359458 176712 359464 176724
rect 355008 176684 359464 176712
rect 355008 176672 355014 176684
rect 359458 176672 359464 176684
rect 359516 176672 359522 176724
rect 362862 176672 362868 176724
rect 362920 176712 362926 176724
rect 363598 176712 363604 176724
rect 362920 176684 363604 176712
rect 362920 176672 362926 176684
rect 363598 176672 363604 176684
rect 363656 176672 363662 176724
rect 368842 176672 368848 176724
rect 368900 176712 368906 176724
rect 371878 176712 371884 176724
rect 368900 176684 371884 176712
rect 368900 176672 368906 176684
rect 371878 176672 371884 176684
rect 371936 176672 371942 176724
rect 380710 176672 380716 176724
rect 380768 176712 380774 176724
rect 381538 176712 381544 176724
rect 380768 176684 381544 176712
rect 380768 176672 380774 176684
rect 381538 176672 381544 176684
rect 381596 176672 381602 176724
rect 384482 176672 384488 176724
rect 384540 176712 384546 176724
rect 385586 176712 385592 176724
rect 384540 176684 385592 176712
rect 384540 176672 384546 176684
rect 385586 176672 385592 176684
rect 385644 176672 385650 176724
rect 327350 176604 327356 176656
rect 327408 176644 327414 176656
rect 327534 176644 327540 176656
rect 327408 176616 327540 176644
rect 327408 176604 327414 176616
rect 327534 176604 327540 176616
rect 327592 176604 327598 176656
rect 357710 176604 357716 176656
rect 357768 176644 357774 176656
rect 357894 176644 357900 176656
rect 357768 176616 357900 176644
rect 357768 176604 357774 176616
rect 357894 176604 357900 176616
rect 357952 176604 357958 176656
rect 309594 175992 309600 176044
rect 309652 176032 309658 176044
rect 394694 176032 394700 176044
rect 309652 176004 394700 176032
rect 309652 175992 309658 176004
rect 394694 175992 394700 176004
rect 394752 175992 394758 176044
rect 125594 175924 125600 175976
rect 125652 175964 125658 175976
rect 223758 175964 223764 175976
rect 125652 175936 223764 175964
rect 125652 175924 125658 175936
rect 223758 175924 223764 175936
rect 223816 175924 223822 175976
rect 275922 175924 275928 175976
rect 275980 175964 275986 175976
rect 316034 175964 316040 175976
rect 275980 175936 316040 175964
rect 275980 175924 275986 175936
rect 316034 175924 316040 175936
rect 316092 175924 316098 175976
rect 390370 175924 390376 175976
rect 390428 175964 390434 175976
rect 579614 175964 579620 175976
rect 390428 175936 579620 175964
rect 390428 175924 390434 175936
rect 579614 175924 579620 175936
rect 579672 175924 579678 175976
rect 340966 175652 340972 175704
rect 341024 175692 341030 175704
rect 341886 175692 341892 175704
rect 341024 175664 341892 175692
rect 341024 175652 341030 175664
rect 341886 175652 341892 175664
rect 341944 175652 341950 175704
rect 375374 175652 375380 175704
rect 375432 175692 375438 175704
rect 376294 175692 376300 175704
rect 375432 175664 376300 175692
rect 375432 175652 375438 175664
rect 376294 175652 376300 175664
rect 376352 175652 376358 175704
rect 194594 175584 194600 175636
rect 194652 175624 194658 175636
rect 194778 175624 194784 175636
rect 194652 175596 194784 175624
rect 194652 175584 194658 175596
rect 194778 175584 194784 175596
rect 194836 175584 194842 175636
rect 200206 175584 200212 175636
rect 200264 175624 200270 175636
rect 201126 175624 201132 175636
rect 200264 175596 201132 175624
rect 200264 175584 200270 175596
rect 201126 175584 201132 175596
rect 201184 175584 201190 175636
rect 207198 175584 207204 175636
rect 207256 175624 207262 175636
rect 207750 175624 207756 175636
rect 207256 175596 207756 175624
rect 207256 175584 207262 175596
rect 207750 175584 207756 175596
rect 207808 175584 207814 175636
rect 215294 175584 215300 175636
rect 215352 175624 215358 175636
rect 215570 175624 215576 175636
rect 215352 175596 215576 175624
rect 215352 175584 215358 175596
rect 215570 175584 215576 175596
rect 215628 175584 215634 175636
rect 218054 175584 218060 175636
rect 218112 175624 218118 175636
rect 218606 175624 218612 175636
rect 218112 175596 218612 175624
rect 218112 175584 218118 175596
rect 218606 175584 218612 175596
rect 218664 175584 218670 175636
rect 229186 175584 229192 175636
rect 229244 175624 229250 175636
rect 230014 175624 230020 175636
rect 229244 175596 230020 175624
rect 229244 175584 229250 175596
rect 230014 175584 230020 175596
rect 230072 175584 230078 175636
rect 230474 175584 230480 175636
rect 230532 175624 230538 175636
rect 230934 175624 230940 175636
rect 230532 175596 230940 175624
rect 230532 175584 230538 175596
rect 230934 175584 230940 175596
rect 230992 175584 230998 175636
rect 233326 175584 233332 175636
rect 233384 175624 233390 175636
rect 234062 175624 234068 175636
rect 233384 175596 234068 175624
rect 233384 175584 233390 175596
rect 234062 175584 234068 175596
rect 234120 175584 234126 175636
rect 241698 175584 241704 175636
rect 241756 175624 241762 175636
rect 242342 175624 242348 175636
rect 241756 175596 242348 175624
rect 241756 175584 241762 175596
rect 242342 175584 242348 175596
rect 242400 175584 242406 175636
rect 242894 175584 242900 175636
rect 242952 175624 242958 175636
rect 243446 175624 243452 175636
rect 242952 175596 243452 175624
rect 242952 175584 242958 175596
rect 243446 175584 243452 175596
rect 243504 175584 243510 175636
rect 253934 175584 253940 175636
rect 253992 175624 253998 175636
rect 254670 175624 254676 175636
rect 253992 175596 254676 175624
rect 253992 175584 253998 175596
rect 254670 175584 254676 175596
rect 254728 175584 254734 175636
rect 255314 175584 255320 175636
rect 255372 175624 255378 175636
rect 256326 175624 256332 175636
rect 255372 175596 256332 175624
rect 255372 175584 255378 175596
rect 256326 175584 256332 175596
rect 256384 175584 256390 175636
rect 259546 175584 259552 175636
rect 259604 175624 259610 175636
rect 260374 175624 260380 175636
rect 259604 175596 260380 175624
rect 259604 175584 259610 175596
rect 260374 175584 260380 175596
rect 260432 175584 260438 175636
rect 263686 175584 263692 175636
rect 263744 175624 263750 175636
rect 264606 175624 264612 175636
rect 263744 175596 264612 175624
rect 263744 175584 263750 175596
rect 264606 175584 264612 175596
rect 264664 175584 264670 175636
rect 267826 175584 267832 175636
rect 267884 175624 267890 175636
rect 268654 175624 268660 175636
rect 267884 175596 268660 175624
rect 267884 175584 267890 175596
rect 268654 175584 268660 175596
rect 268712 175584 268718 175636
rect 269114 175584 269120 175636
rect 269172 175624 269178 175636
rect 269758 175624 269764 175636
rect 269172 175596 269764 175624
rect 269172 175584 269178 175596
rect 269758 175584 269764 175596
rect 269816 175584 269822 175636
rect 287054 175584 287060 175636
rect 287112 175624 287118 175636
rect 287790 175624 287796 175636
rect 287112 175596 287796 175624
rect 287112 175584 287118 175596
rect 287790 175584 287796 175596
rect 287848 175584 287854 175636
rect 302326 175584 302332 175636
rect 302384 175624 302390 175636
rect 303246 175624 303252 175636
rect 302384 175596 303252 175624
rect 302384 175584 302390 175596
rect 303246 175584 303252 175596
rect 303304 175584 303310 175636
rect 305178 175584 305184 175636
rect 305236 175624 305242 175636
rect 305822 175624 305828 175636
rect 305236 175596 305828 175624
rect 305236 175584 305242 175596
rect 305822 175584 305828 175596
rect 305880 175584 305886 175636
rect 310514 175584 310520 175636
rect 310572 175624 310578 175636
rect 311342 175624 311348 175636
rect 310572 175596 311348 175624
rect 310572 175584 310578 175596
rect 311342 175584 311348 175596
rect 311400 175584 311406 175636
rect 311894 175584 311900 175636
rect 311952 175624 311958 175636
rect 312446 175624 312452 175636
rect 311952 175596 312452 175624
rect 311952 175584 311958 175596
rect 312446 175584 312452 175596
rect 312504 175584 312510 175636
rect 340874 175584 340880 175636
rect 340932 175624 340938 175636
rect 341334 175624 341340 175636
rect 340932 175596 341340 175624
rect 340932 175584 340938 175596
rect 341334 175584 341340 175596
rect 341392 175584 341398 175636
rect 342254 175584 342260 175636
rect 342312 175624 342318 175636
rect 342806 175624 342812 175636
rect 342312 175596 342812 175624
rect 342312 175584 342318 175596
rect 342806 175584 342812 175596
rect 342864 175584 342870 175636
rect 343634 175584 343640 175636
rect 343692 175624 343698 175636
rect 344462 175624 344468 175636
rect 343692 175596 344468 175624
rect 343692 175584 343698 175596
rect 344462 175584 344468 175596
rect 344520 175584 344526 175636
rect 345014 175584 345020 175636
rect 345072 175624 345078 175636
rect 345934 175624 345940 175636
rect 345072 175596 345940 175624
rect 345072 175584 345078 175596
rect 345934 175584 345940 175596
rect 345992 175584 345998 175636
rect 347774 175584 347780 175636
rect 347832 175624 347838 175636
rect 348510 175624 348516 175636
rect 347832 175596 348516 175624
rect 347832 175584 347838 175596
rect 348510 175584 348516 175596
rect 348568 175584 348574 175636
rect 349154 175584 349160 175636
rect 349212 175624 349218 175636
rect 350166 175624 350172 175636
rect 349212 175596 350172 175624
rect 349212 175584 349218 175596
rect 350166 175584 350172 175596
rect 350224 175584 350230 175636
rect 362954 175584 362960 175636
rect 363012 175624 363018 175636
rect 363414 175624 363420 175636
rect 363012 175596 363420 175624
rect 363012 175584 363018 175596
rect 363414 175584 363420 175596
rect 363472 175584 363478 175636
rect 375466 175584 375472 175636
rect 375524 175624 375530 175636
rect 375926 175624 375932 175636
rect 375524 175596 375932 175624
rect 375524 175584 375530 175596
rect 375926 175584 375932 175596
rect 375984 175584 375990 175636
rect 249794 175516 249800 175568
rect 249852 175556 249858 175568
rect 250070 175556 250076 175568
rect 249852 175528 250076 175556
rect 249852 175516 249858 175528
rect 250070 175516 250076 175528
rect 250128 175516 250134 175568
rect 288434 175516 288440 175568
rect 288492 175556 288498 175568
rect 289262 175556 289268 175568
rect 288492 175528 289268 175556
rect 288492 175516 288498 175528
rect 289262 175516 289268 175528
rect 289320 175516 289326 175568
rect 313366 175516 313372 175568
rect 313424 175556 313430 175568
rect 313918 175556 313924 175568
rect 313424 175528 313924 175556
rect 313424 175516 313430 175528
rect 313918 175516 313924 175528
rect 313976 175516 313982 175568
rect 317506 175516 317512 175568
rect 317564 175556 317570 175568
rect 318150 175556 318156 175568
rect 317564 175528 318156 175556
rect 317564 175516 317570 175528
rect 318150 175516 318156 175528
rect 318208 175516 318214 175568
rect 284294 175448 284300 175500
rect 284352 175488 284358 175500
rect 284662 175488 284668 175500
rect 284352 175460 284668 175488
rect 284352 175448 284358 175460
rect 284662 175448 284668 175460
rect 284720 175448 284726 175500
rect 339494 175448 339500 175500
rect 339552 175488 339558 175500
rect 339862 175488 339868 175500
rect 339552 175460 339868 175488
rect 339552 175448 339558 175460
rect 339862 175448 339868 175460
rect 339920 175448 339926 175500
rect 373994 175448 374000 175500
rect 374052 175488 374058 175500
rect 374822 175488 374828 175500
rect 374052 175460 374828 175488
rect 374052 175448 374058 175460
rect 374822 175448 374828 175460
rect 374880 175448 374886 175500
rect 160094 174564 160100 174616
rect 160152 174604 160158 174616
rect 207014 174604 207020 174616
rect 160152 174576 207020 174604
rect 160152 174564 160158 174576
rect 207014 174564 207020 174576
rect 207072 174564 207078 174616
rect 348418 174564 348424 174616
rect 348476 174604 348482 174616
rect 483014 174604 483020 174616
rect 348476 174576 483020 174604
rect 348476 174564 348482 174576
rect 483014 174564 483020 174576
rect 483072 174564 483078 174616
rect 155218 174496 155224 174548
rect 155276 174536 155282 174548
rect 202874 174536 202880 174548
rect 155276 174508 202880 174536
rect 155276 174496 155282 174508
rect 202874 174496 202880 174508
rect 202932 174496 202938 174548
rect 283650 174496 283656 174548
rect 283708 174536 283714 174548
rect 333974 174536 333980 174548
rect 283708 174508 333980 174536
rect 283708 174496 283714 174508
rect 333974 174496 333980 174508
rect 334032 174496 334038 174548
rect 387702 174496 387708 174548
rect 387760 174536 387766 174548
rect 571978 174536 571984 174548
rect 387760 174508 571984 174536
rect 387760 174496 387766 174508
rect 571978 174496 571984 174508
rect 572036 174496 572042 174548
rect 258258 174088 258264 174140
rect 258316 174128 258322 174140
rect 258902 174128 258908 174140
rect 258316 174100 258908 174128
rect 258316 174088 258322 174100
rect 258902 174088 258908 174100
rect 258960 174088 258966 174140
rect 236086 173952 236092 174004
rect 236144 173992 236150 174004
rect 236270 173992 236276 174004
rect 236144 173964 236276 173992
rect 236144 173952 236150 173964
rect 236270 173952 236276 173964
rect 236328 173952 236334 174004
rect 346394 173816 346400 173868
rect 346452 173856 346458 173868
rect 347038 173856 347044 173868
rect 346452 173828 347044 173856
rect 346452 173816 346458 173828
rect 347038 173816 347044 173828
rect 347096 173816 347102 173868
rect 164234 173204 164240 173256
rect 164292 173244 164298 173256
rect 208394 173244 208400 173256
rect 164292 173216 208400 173244
rect 164292 173204 164298 173216
rect 208394 173204 208400 173216
rect 208452 173204 208458 173256
rect 333330 173204 333336 173256
rect 333388 173244 333394 173256
rect 448514 173244 448520 173256
rect 333388 173216 448520 173244
rect 333388 173204 333394 173216
rect 448514 173204 448520 173216
rect 448572 173204 448578 173256
rect 158714 173136 158720 173188
rect 158772 173176 158778 173188
rect 205634 173176 205640 173188
rect 158772 173148 205640 173176
rect 158772 173136 158778 173148
rect 205634 173136 205640 173148
rect 205692 173136 205698 173188
rect 279142 173136 279148 173188
rect 279200 173176 279206 173188
rect 324406 173176 324412 173188
rect 279200 173148 324412 173176
rect 279200 173136 279206 173148
rect 324406 173136 324412 173148
rect 324464 173136 324470 173188
rect 351730 173136 351736 173188
rect 351788 173176 351794 173188
rect 489914 173176 489920 173188
rect 351788 173148 489920 173176
rect 351788 173136 351794 173148
rect 489914 173136 489920 173148
rect 489972 173136 489978 173188
rect 209958 171980 209964 172032
rect 210016 172020 210022 172032
rect 226334 172020 226340 172032
rect 210016 171992 226340 172020
rect 210016 171980 210022 171992
rect 226334 171980 226340 171992
rect 226392 171980 226398 172032
rect 168374 171844 168380 171896
rect 168432 171884 168438 171896
rect 209774 171884 209780 171896
rect 168432 171856 209780 171884
rect 168432 171844 168438 171856
rect 209774 171844 209780 171856
rect 209832 171844 209838 171896
rect 314746 171844 314752 171896
rect 314804 171884 314810 171896
rect 407114 171884 407120 171896
rect 314804 171856 407120 171884
rect 314804 171844 314810 171856
rect 407114 171844 407120 171856
rect 407172 171844 407178 171896
rect 142798 171776 142804 171828
rect 142856 171816 142862 171828
rect 197998 171816 198004 171828
rect 142856 171788 198004 171816
rect 142856 171776 142862 171788
rect 197998 171776 198004 171788
rect 198056 171776 198062 171828
rect 248506 171776 248512 171828
rect 248564 171816 248570 171828
rect 248966 171816 248972 171828
rect 248564 171788 248972 171816
rect 248564 171776 248570 171788
rect 248966 171776 248972 171788
rect 249024 171776 249030 171828
rect 273254 171776 273260 171828
rect 273312 171816 273318 171828
rect 273806 171816 273812 171828
rect 273312 171788 273812 171816
rect 273312 171776 273318 171788
rect 273806 171776 273812 171788
rect 273864 171776 273870 171828
rect 280154 171776 280160 171828
rect 280212 171816 280218 171828
rect 280430 171816 280436 171828
rect 280212 171788 280436 171816
rect 280212 171776 280218 171788
rect 280430 171776 280436 171788
rect 280488 171776 280494 171828
rect 292574 171776 292580 171828
rect 292632 171816 292638 171828
rect 293310 171816 293316 171828
rect 292632 171788 293316 171816
rect 292632 171776 292638 171788
rect 293310 171776 293316 171788
rect 293368 171776 293374 171828
rect 298094 171776 298100 171828
rect 298152 171816 298158 171828
rect 299014 171816 299020 171828
rect 298152 171788 299020 171816
rect 298152 171776 298158 171788
rect 299014 171776 299020 171788
rect 299072 171776 299078 171828
rect 299474 171776 299480 171828
rect 299532 171816 299538 171828
rect 300118 171816 300124 171828
rect 299532 171788 300124 171816
rect 299532 171776 299538 171788
rect 300118 171776 300124 171788
rect 300176 171776 300182 171828
rect 322934 171776 322940 171828
rect 322992 171816 322998 171828
rect 323854 171816 323860 171828
rect 322992 171788 323860 171816
rect 322992 171776 322998 171788
rect 323854 171776 323860 171788
rect 323912 171776 323918 171828
rect 327166 171776 327172 171828
rect 327224 171816 327230 171828
rect 327902 171816 327908 171828
rect 327224 171788 327908 171816
rect 327224 171776 327230 171788
rect 327902 171776 327908 171788
rect 327960 171776 327966 171828
rect 353294 171776 353300 171828
rect 353352 171816 353358 171828
rect 353662 171816 353668 171828
rect 353352 171788 353668 171816
rect 353352 171776 353358 171788
rect 353662 171776 353668 171788
rect 353720 171776 353726 171828
rect 356146 171776 356152 171828
rect 356204 171816 356210 171828
rect 356790 171816 356796 171828
rect 356204 171788 356796 171816
rect 356204 171776 356210 171788
rect 356790 171776 356796 171788
rect 356848 171776 356854 171828
rect 357434 171776 357440 171828
rect 357492 171816 357498 171828
rect 358262 171816 358268 171828
rect 357492 171788 358268 171816
rect 357492 171776 357498 171788
rect 358262 171776 358268 171788
rect 358320 171776 358326 171828
rect 494054 171816 494060 171828
rect 360166 171788 494060 171816
rect 353386 171708 353392 171760
rect 353444 171748 353450 171760
rect 354214 171748 354220 171760
rect 353444 171720 354220 171748
rect 353444 171708 353450 171720
rect 354214 171708 354220 171720
rect 354272 171708 354278 171760
rect 353202 171640 353208 171692
rect 353260 171680 353266 171692
rect 360166 171680 360194 171788
rect 494054 171776 494060 171788
rect 494112 171776 494118 171828
rect 379514 171708 379520 171760
rect 379572 171748 379578 171760
rect 379974 171748 379980 171760
rect 379572 171720 379980 171748
rect 379572 171708 379578 171720
rect 379974 171708 379980 171720
rect 380032 171708 380038 171760
rect 380894 171708 380900 171760
rect 380952 171748 380958 171760
rect 381446 171748 381452 171760
rect 380952 171720 381452 171748
rect 380952 171708 380958 171720
rect 381446 171708 381452 171720
rect 381504 171708 381510 171760
rect 385034 171708 385040 171760
rect 385092 171748 385098 171760
rect 385678 171748 385684 171760
rect 385092 171720 385684 171748
rect 385092 171708 385098 171720
rect 385678 171708 385684 171720
rect 385736 171708 385742 171760
rect 387794 171708 387800 171760
rect 387852 171748 387858 171760
rect 388254 171748 388260 171760
rect 387852 171720 388260 171748
rect 387852 171708 387858 171720
rect 388254 171708 388260 171720
rect 388312 171708 388318 171760
rect 353260 171652 360194 171680
rect 353260 171640 353266 171652
rect 383654 171640 383660 171692
rect 383712 171680 383718 171692
rect 384574 171680 384580 171692
rect 383712 171652 384580 171680
rect 383712 171640 383718 171652
rect 384574 171640 384580 171652
rect 384632 171640 384638 171692
rect 204254 171232 204260 171284
rect 204312 171272 204318 171284
rect 204806 171272 204812 171284
rect 204312 171244 204812 171272
rect 204312 171232 204318 171244
rect 204806 171232 204812 171244
rect 204864 171232 204870 171284
rect 321646 171096 321652 171148
rect 321704 171136 321710 171148
rect 322198 171136 322204 171148
rect 321704 171108 322204 171136
rect 321704 171096 321710 171108
rect 322198 171096 322204 171108
rect 322256 171096 322262 171148
rect 329926 171096 329932 171148
rect 329984 171136 329990 171148
rect 330478 171136 330484 171148
rect 329984 171108 330484 171136
rect 329984 171096 329990 171108
rect 330478 171096 330484 171108
rect 330536 171096 330542 171148
rect 186314 170416 186320 170468
rect 186372 170456 186378 170468
rect 218146 170456 218152 170468
rect 186372 170428 218152 170456
rect 186372 170416 186378 170428
rect 218146 170416 218152 170428
rect 218204 170416 218210 170468
rect 143534 170348 143540 170400
rect 143592 170388 143598 170400
rect 198918 170388 198924 170400
rect 143592 170360 198924 170388
rect 143592 170348 143598 170360
rect 198918 170348 198924 170360
rect 198976 170348 198982 170400
rect 292758 170348 292764 170400
rect 292816 170388 292822 170400
rect 356054 170388 356060 170400
rect 292816 170360 356060 170388
rect 292816 170348 292822 170360
rect 356054 170348 356060 170360
rect 356112 170348 356118 170400
rect 356330 170348 356336 170400
rect 356388 170388 356394 170400
rect 500954 170388 500960 170400
rect 356388 170360 500960 170388
rect 356388 170348 356394 170360
rect 500954 170348 500960 170360
rect 501012 170348 501018 170400
rect 190454 169056 190460 169108
rect 190512 169096 190518 169108
rect 219618 169096 219624 169108
rect 190512 169068 219624 169096
rect 190512 169056 190518 169068
rect 219618 169056 219624 169068
rect 219676 169056 219682 169108
rect 337654 169056 337660 169108
rect 337712 169096 337718 169108
rect 459554 169096 459560 169108
rect 337712 169068 459560 169096
rect 337712 169056 337718 169068
rect 459554 169056 459560 169068
rect 459612 169056 459618 169108
rect 146294 168988 146300 169040
rect 146352 169028 146358 169040
rect 200574 169028 200580 169040
rect 146352 169000 200580 169028
rect 146352 168988 146358 169000
rect 200574 168988 200580 169000
rect 200632 168988 200638 169040
rect 298186 168988 298192 169040
rect 298244 169028 298250 169040
rect 298370 169028 298376 169040
rect 298244 169000 298376 169028
rect 298244 168988 298250 169000
rect 298370 168988 298376 169000
rect 298428 168988 298434 169040
rect 358906 168988 358912 169040
rect 358964 169028 358970 169040
rect 507854 169028 507860 169040
rect 358964 169000 507860 169028
rect 358964 168988 358970 169000
rect 507854 168988 507860 169000
rect 507912 168988 507918 169040
rect 150434 167628 150440 167680
rect 150492 167668 150498 167680
rect 202138 167668 202144 167680
rect 150492 167640 202144 167668
rect 150492 167628 150498 167640
rect 202138 167628 202144 167640
rect 202196 167628 202202 167680
rect 361850 167628 361856 167680
rect 361908 167668 361914 167680
rect 514754 167668 514760 167680
rect 361908 167640 514760 167668
rect 361908 167628 361914 167640
rect 514754 167628 514760 167640
rect 514812 167628 514818 167680
rect 276106 167016 276112 167068
rect 276164 167056 276170 167068
rect 276934 167056 276940 167068
rect 276164 167028 276940 167056
rect 276164 167016 276170 167028
rect 276934 167016 276940 167028
rect 276992 167016 276998 167068
rect 554038 166948 554044 167000
rect 554096 166988 554102 167000
rect 580166 166988 580172 167000
rect 554096 166960 580172 166988
rect 554096 166948 554102 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 297542 166336 297548 166388
rect 297600 166376 297606 166388
rect 367186 166376 367192 166388
rect 297600 166348 367192 166376
rect 297600 166336 297606 166348
rect 367186 166336 367192 166348
rect 367244 166336 367250 166388
rect 157334 166268 157340 166320
rect 157392 166308 157398 166320
rect 205174 166308 205180 166320
rect 157392 166280 205180 166308
rect 157392 166268 157398 166280
rect 205174 166268 205180 166280
rect 205232 166268 205238 166320
rect 366450 166268 366456 166320
rect 366508 166308 366514 166320
rect 525794 166308 525800 166320
rect 366508 166280 525800 166308
rect 366508 166268 366514 166280
rect 525794 166268 525800 166280
rect 525852 166268 525858 166320
rect 311986 164908 311992 164960
rect 312044 164948 312050 164960
rect 400214 164948 400220 164960
rect 312044 164920 400220 164948
rect 312044 164908 312050 164920
rect 400214 164908 400220 164920
rect 400272 164908 400278 164960
rect 161474 164840 161480 164892
rect 161532 164880 161538 164892
rect 207290 164880 207296 164892
rect 161532 164852 207296 164880
rect 161532 164840 161538 164852
rect 207290 164840 207296 164852
rect 207348 164840 207354 164892
rect 368474 164840 368480 164892
rect 368532 164880 368538 164892
rect 529934 164880 529940 164892
rect 368532 164852 529940 164880
rect 368532 164840 368538 164852
rect 529934 164840 529940 164852
rect 529992 164840 529998 164892
rect 3326 164160 3332 164212
rect 3384 164200 3390 164212
rect 14458 164200 14464 164212
rect 3384 164172 14464 164200
rect 3384 164160 3390 164172
rect 14458 164160 14464 164172
rect 14516 164160 14522 164212
rect 308306 163548 308312 163600
rect 308364 163588 308370 163600
rect 391934 163588 391940 163600
rect 308364 163560 391940 163588
rect 308364 163548 308370 163560
rect 391934 163548 391940 163560
rect 391992 163548 391998 163600
rect 165614 163480 165620 163532
rect 165672 163520 165678 163532
rect 208486 163520 208492 163532
rect 165672 163492 208492 163520
rect 165672 163480 165678 163492
rect 208486 163480 208492 163492
rect 208544 163480 208550 163532
rect 372798 163480 372804 163532
rect 372856 163520 372862 163532
rect 539594 163520 539600 163532
rect 372856 163492 539600 163520
rect 372856 163480 372862 163492
rect 539594 163480 539600 163492
rect 539652 163480 539658 163532
rect 319070 162188 319076 162240
rect 319128 162228 319134 162240
rect 416774 162228 416780 162240
rect 319128 162200 416780 162228
rect 319128 162188 319134 162200
rect 416774 162188 416780 162200
rect 416832 162188 416838 162240
rect 172514 162120 172520 162172
rect 172572 162160 172578 162172
rect 211890 162160 211896 162172
rect 172572 162132 211896 162160
rect 172572 162120 172578 162132
rect 211890 162120 211896 162132
rect 211948 162120 211954 162172
rect 374178 162120 374184 162172
rect 374236 162160 374242 162172
rect 543734 162160 543740 162172
rect 374236 162132 543740 162160
rect 374236 162120 374242 162132
rect 543734 162120 543740 162132
rect 543792 162120 543798 162172
rect 316218 160760 316224 160812
rect 316276 160800 316282 160812
rect 411254 160800 411260 160812
rect 316276 160772 411260 160800
rect 316276 160760 316282 160772
rect 411254 160760 411260 160772
rect 411312 160760 411318 160812
rect 176746 160692 176752 160744
rect 176804 160732 176810 160744
rect 212718 160732 212724 160744
rect 176804 160704 212724 160732
rect 176804 160692 176810 160704
rect 212718 160692 212724 160704
rect 212776 160692 212782 160744
rect 375466 160692 375472 160744
rect 375524 160732 375530 160744
rect 547874 160732 547880 160744
rect 375524 160704 547880 160732
rect 375524 160692 375530 160704
rect 547874 160692 547880 160704
rect 547932 160692 547938 160744
rect 328454 159400 328460 159452
rect 328512 159440 328518 159452
rect 438854 159440 438860 159452
rect 328512 159412 438860 159440
rect 328512 159400 328518 159412
rect 438854 159400 438860 159412
rect 438912 159400 438918 159452
rect 179414 159332 179420 159384
rect 179472 159372 179478 159384
rect 215478 159372 215484 159384
rect 179472 159344 215484 159372
rect 179472 159332 179478 159344
rect 215478 159332 215484 159344
rect 215536 159332 215542 159384
rect 378410 159332 378416 159384
rect 378468 159372 378474 159384
rect 554774 159372 554780 159384
rect 378468 159344 554780 159372
rect 378468 159332 378474 159344
rect 554774 159332 554780 159344
rect 554832 159332 554838 159384
rect 327258 158040 327264 158092
rect 327316 158080 327322 158092
rect 434714 158080 434720 158092
rect 327316 158052 434720 158080
rect 327316 158040 327322 158052
rect 434714 158040 434720 158052
rect 434772 158040 434778 158092
rect 183554 157972 183560 158024
rect 183612 158012 183618 158024
rect 216766 158012 216772 158024
rect 183612 157984 216772 158012
rect 183612 157972 183618 157984
rect 216766 157972 216772 157984
rect 216824 157972 216830 158024
rect 381538 157972 381544 158024
rect 381596 158012 381602 158024
rect 557534 158012 557540 158024
rect 381596 157984 557540 158012
rect 381596 157972 381602 157984
rect 557534 157972 557540 157984
rect 557592 157972 557598 158024
rect 314654 156680 314660 156732
rect 314712 156720 314718 156732
rect 407206 156720 407212 156732
rect 314712 156692 407212 156720
rect 314712 156680 314718 156692
rect 407206 156680 407212 156692
rect 407264 156680 407270 156732
rect 129734 156612 129740 156664
rect 129792 156652 129798 156664
rect 192478 156652 192484 156664
rect 129792 156624 192484 156652
rect 129792 156612 129798 156624
rect 192478 156612 192484 156624
rect 192536 156612 192542 156664
rect 382182 156612 382188 156664
rect 382240 156652 382246 156664
rect 561674 156652 561680 156664
rect 382240 156624 561680 156652
rect 382240 156612 382246 156624
rect 561674 156612 561680 156624
rect 561732 156612 561738 156664
rect 313458 155252 313464 155304
rect 313516 155292 313522 155304
rect 404354 155292 404360 155304
rect 313516 155264 404360 155292
rect 313516 155252 313522 155264
rect 404354 155252 404360 155264
rect 404412 155252 404418 155304
rect 137278 155184 137284 155236
rect 137336 155224 137342 155236
rect 194686 155224 194692 155236
rect 137336 155196 194692 155224
rect 137336 155184 137342 155196
rect 194686 155184 194692 155196
rect 194744 155184 194750 155236
rect 383746 155184 383752 155236
rect 383804 155224 383810 155236
rect 564434 155224 564440 155236
rect 383804 155196 564440 155224
rect 383804 155184 383810 155196
rect 564434 155184 564440 155196
rect 564492 155184 564498 155236
rect 309226 153892 309232 153944
rect 309284 153932 309290 153944
rect 396074 153932 396080 153944
rect 309284 153904 396080 153932
rect 309284 153892 309290 153904
rect 396074 153892 396080 153904
rect 396132 153892 396138 153944
rect 140038 153824 140044 153876
rect 140096 153864 140102 153876
rect 196066 153864 196072 153876
rect 140096 153836 196072 153864
rect 140096 153824 140102 153836
rect 196066 153824 196072 153836
rect 196124 153824 196130 153876
rect 385126 153824 385132 153876
rect 385184 153864 385190 153876
rect 568574 153864 568580 153876
rect 385184 153836 568580 153864
rect 385184 153824 385190 153836
rect 568574 153824 568580 153836
rect 568632 153824 568638 153876
rect 394510 153144 394516 153196
rect 394568 153184 394574 153196
rect 580166 153184 580172 153196
rect 394568 153156 580172 153184
rect 394568 153144 394574 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 148318 152464 148324 152516
rect 148376 152504 148382 152516
rect 199010 152504 199016 152516
rect 148376 152476 199016 152504
rect 148376 152464 148382 152476
rect 199010 152464 199016 152476
rect 199068 152464 199074 152516
rect 306466 152464 306472 152516
rect 306524 152504 306530 152516
rect 389174 152504 389180 152516
rect 306524 152476 389180 152504
rect 306524 152464 306530 152476
rect 389174 152464 389180 152476
rect 389232 152464 389238 152516
rect 152458 151036 152464 151088
rect 152516 151076 152522 151088
rect 200206 151076 200212 151088
rect 152516 151048 200212 151076
rect 152516 151036 152522 151048
rect 200206 151036 200212 151048
rect 200264 151036 200270 151088
rect 386598 151036 386604 151088
rect 386656 151076 386662 151088
rect 572806 151076 572812 151088
rect 386656 151048 572812 151076
rect 386656 151036 386662 151048
rect 572806 151036 572812 151048
rect 572864 151036 572870 151088
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 190178 150396 190184 150408
rect 3384 150368 190184 150396
rect 3384 150356 3390 150368
rect 190178 150356 190184 150368
rect 190236 150356 190242 150408
rect 310790 149744 310796 149796
rect 310848 149784 310854 149796
rect 398834 149784 398840 149796
rect 310848 149756 398840 149784
rect 310848 149744 310854 149756
rect 398834 149744 398840 149756
rect 398892 149744 398898 149796
rect 379606 149676 379612 149728
rect 379664 149716 379670 149728
rect 556154 149716 556160 149728
rect 379664 149688 556160 149716
rect 379664 149676 379670 149688
rect 556154 149676 556160 149688
rect 556212 149676 556218 149728
rect 321738 148384 321744 148436
rect 321796 148424 321802 148436
rect 423674 148424 423680 148436
rect 321796 148396 423680 148424
rect 321796 148384 321802 148396
rect 423674 148384 423680 148396
rect 423732 148384 423738 148436
rect 156598 148316 156604 148368
rect 156656 148356 156662 148368
rect 204346 148356 204352 148368
rect 156656 148328 204352 148356
rect 156656 148316 156662 148328
rect 204346 148316 204352 148328
rect 204404 148316 204410 148368
rect 387978 148316 387984 148368
rect 388036 148356 388042 148368
rect 574738 148356 574744 148368
rect 388036 148328 574744 148356
rect 388036 148316 388042 148328
rect 574738 148316 574744 148328
rect 574796 148316 574802 148368
rect 324498 146956 324504 147008
rect 324556 146996 324562 147008
rect 430574 146996 430580 147008
rect 324556 146968 430580 146996
rect 324556 146956 324562 146968
rect 430574 146956 430580 146968
rect 430632 146956 430638 147008
rect 367278 146888 367284 146940
rect 367336 146928 367342 146940
rect 528554 146928 528560 146940
rect 367336 146900 528560 146928
rect 367336 146888 367342 146900
rect 528554 146888 528560 146900
rect 528612 146888 528618 146940
rect 329834 145528 329840 145580
rect 329892 145568 329898 145580
rect 440326 145568 440332 145580
rect 329892 145540 440332 145568
rect 329892 145528 329898 145540
rect 440326 145528 440332 145540
rect 440384 145528 440390 145580
rect 335998 144168 336004 144220
rect 336056 144208 336062 144220
rect 448606 144208 448612 144220
rect 336056 144180 448612 144208
rect 336056 144168 336062 144180
rect 448606 144168 448612 144180
rect 448664 144168 448670 144220
rect 338850 142808 338856 142860
rect 338908 142848 338914 142860
rect 458174 142848 458180 142860
rect 338908 142820 458180 142848
rect 338908 142808 338914 142820
rect 458174 142808 458180 142820
rect 458232 142808 458238 142860
rect 347774 141380 347780 141432
rect 347832 141420 347838 141432
rect 484394 141420 484400 141432
rect 347832 141392 484400 141420
rect 347832 141380 347838 141392
rect 484394 141380 484400 141392
rect 484452 141380 484458 141432
rect 353478 140020 353484 140072
rect 353536 140060 353542 140072
rect 495434 140060 495440 140072
rect 353536 140032 495440 140060
rect 353536 140020 353542 140032
rect 495434 140020 495440 140032
rect 495492 140020 495498 140072
rect 399478 139340 399484 139392
rect 399536 139380 399542 139392
rect 579890 139380 579896 139392
rect 399536 139352 579896 139380
rect 399536 139340 399542 139352
rect 579890 139340 579896 139352
rect 579948 139340 579954 139392
rect 3050 137912 3056 137964
rect 3108 137952 3114 137964
rect 189994 137952 190000 137964
rect 3108 137924 190000 137952
rect 3108 137912 3114 137924
rect 189994 137912 190000 137924
rect 190052 137912 190058 137964
rect 356238 137232 356244 137284
rect 356296 137272 356302 137284
rect 502334 137272 502340 137284
rect 356296 137244 502340 137272
rect 356296 137232 356302 137244
rect 502334 137232 502340 137244
rect 502392 137232 502398 137284
rect 357526 135872 357532 135924
rect 357584 135912 357590 135924
rect 506474 135912 506480 135924
rect 357584 135884 506480 135912
rect 357584 135872 357590 135884
rect 506474 135872 506480 135884
rect 506532 135872 506538 135924
rect 360378 134512 360384 134564
rect 360436 134552 360442 134564
rect 513374 134552 513380 134564
rect 360436 134524 513380 134552
rect 360436 134512 360442 134524
rect 513374 134512 513380 134524
rect 513432 134512 513438 134564
rect 363598 133152 363604 133204
rect 363656 133192 363662 133204
rect 516134 133192 516140 133204
rect 363656 133164 516140 133192
rect 363656 133152 363662 133164
rect 516134 133152 516140 133164
rect 516192 133152 516198 133204
rect 364334 131724 364340 131776
rect 364392 131764 364398 131776
rect 520274 131764 520280 131776
rect 364392 131736 520280 131764
rect 364392 131724 364398 131736
rect 520274 131724 520280 131736
rect 520332 131724 520338 131776
rect 374638 130364 374644 130416
rect 374696 130404 374702 130416
rect 540974 130404 540980 130416
rect 374696 130376 540980 130404
rect 374696 130364 374702 130376
rect 540974 130364 540980 130376
rect 541032 130364 541038 130416
rect 305270 129004 305276 129056
rect 305328 129044 305334 129056
rect 385126 129044 385132 129056
rect 305328 129016 385132 129044
rect 305328 129004 305334 129016
rect 385126 129004 385132 129016
rect 385184 129004 385190 129056
rect 385678 129004 385684 129056
rect 385736 129044 385742 129056
rect 565814 129044 565820 129056
rect 385736 129016 565820 129044
rect 385736 129004 385742 129016
rect 565814 129004 565820 129016
rect 565872 129004 565878 129056
rect 312538 127576 312544 127628
rect 312596 127616 312602 127628
rect 376846 127616 376852 127628
rect 312596 127588 376852 127616
rect 312596 127576 312602 127588
rect 376846 127576 376852 127588
rect 376904 127576 376910 127628
rect 380986 127576 380992 127628
rect 381044 127616 381050 127628
rect 558914 127616 558920 127628
rect 381044 127588 558920 127616
rect 381044 127576 381050 127588
rect 558914 127576 558920 127588
rect 558972 127576 558978 127628
rect 551278 126896 551284 126948
rect 551336 126936 551342 126948
rect 579982 126936 579988 126948
rect 551336 126908 579988 126936
rect 551336 126896 551342 126908
rect 579982 126896 579988 126908
rect 580040 126896 580046 126948
rect 376938 126216 376944 126268
rect 376996 126256 377002 126268
rect 550634 126256 550640 126268
rect 376996 126228 550640 126256
rect 376996 126216 377002 126228
rect 550634 126216 550640 126228
rect 550692 126216 550698 126268
rect 325694 124856 325700 124908
rect 325752 124896 325758 124908
rect 432046 124896 432052 124908
rect 325752 124868 432052 124896
rect 325752 124856 325758 124868
rect 432046 124856 432052 124868
rect 432104 124856 432110 124908
rect 280430 123428 280436 123480
rect 280488 123468 280494 123480
rect 329834 123468 329840 123480
rect 280488 123440 329840 123468
rect 280488 123428 280494 123440
rect 329834 123428 329840 123440
rect 329892 123428 329898 123480
rect 330018 123428 330024 123480
rect 330076 123468 330082 123480
rect 441614 123468 441620 123480
rect 330076 123440 441620 123468
rect 330076 123428 330082 123440
rect 441614 123428 441620 123440
rect 441672 123428 441678 123480
rect 331398 122068 331404 122120
rect 331456 122108 331462 122120
rect 445754 122108 445760 122120
rect 331456 122080 445760 122108
rect 331456 122068 331462 122080
rect 445754 122068 445760 122080
rect 445812 122068 445818 122120
rect 334158 120708 334164 120760
rect 334216 120748 334222 120760
rect 452654 120748 452660 120760
rect 334216 120720 452660 120748
rect 334216 120708 334222 120720
rect 452654 120708 452660 120720
rect 452712 120708 452718 120760
rect 339586 119348 339592 119400
rect 339644 119388 339650 119400
rect 463694 119388 463700 119400
rect 339644 119360 463700 119388
rect 339644 119348 339650 119360
rect 463694 119348 463700 119360
rect 463752 119348 463758 119400
rect 343818 117920 343824 117972
rect 343876 117960 343882 117972
rect 473354 117960 473360 117972
rect 343876 117932 473360 117960
rect 343876 117920 343882 117932
rect 473354 117920 473360 117932
rect 473412 117920 473418 117972
rect 347866 116628 347872 116680
rect 347924 116668 347930 116680
rect 347924 116640 354674 116668
rect 347924 116628 347930 116640
rect 288618 116560 288624 116612
rect 288676 116600 288682 116612
rect 347774 116600 347780 116612
rect 288676 116572 347780 116600
rect 288676 116560 288682 116572
rect 347774 116560 347780 116572
rect 347832 116560 347838 116612
rect 354646 116600 354674 116640
rect 481634 116600 481640 116612
rect 354646 116572 481640 116600
rect 481634 116560 481640 116572
rect 481692 116560 481698 116612
rect 350534 115200 350540 115252
rect 350592 115240 350598 115252
rect 490006 115240 490012 115252
rect 350592 115212 490012 115240
rect 350592 115200 350598 115212
rect 490006 115200 490012 115212
rect 490064 115200 490070 115252
rect 354674 113772 354680 113824
rect 354732 113812 354738 113824
rect 499574 113812 499580 113824
rect 354732 113784 499580 113812
rect 354732 113772 354738 113784
rect 499574 113772 499580 113784
rect 499632 113772 499638 113824
rect 394418 113092 394424 113144
rect 394476 113132 394482 113144
rect 580166 113132 580172 113144
rect 394476 113104 580172 113132
rect 394476 113092 394482 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 361574 111052 361580 111104
rect 361632 111092 361638 111104
rect 514846 111092 514852 111104
rect 361632 111064 514852 111092
rect 361632 111052 361638 111064
rect 514846 111052 514852 111064
rect 514904 111052 514910 111104
rect 3326 110848 3332 110900
rect 3384 110888 3390 110900
rect 7558 110888 7564 110900
rect 3384 110860 7564 110888
rect 3384 110848 3390 110860
rect 7558 110848 7564 110860
rect 7616 110848 7622 110900
rect 365806 109692 365812 109744
rect 365864 109732 365870 109744
rect 524414 109732 524420 109744
rect 365864 109704 524420 109732
rect 365864 109692 365870 109704
rect 524414 109692 524420 109704
rect 524472 109692 524478 109744
rect 370130 108264 370136 108316
rect 370188 108304 370194 108316
rect 535454 108304 535460 108316
rect 370188 108276 535460 108304
rect 370188 108264 370194 108276
rect 535454 108264 535460 108276
rect 535512 108264 535518 108316
rect 372614 106904 372620 106956
rect 372672 106944 372678 106956
rect 539686 106944 539692 106956
rect 372672 106916 539692 106944
rect 372672 106904 372678 106916
rect 539686 106904 539692 106916
rect 539744 106904 539750 106956
rect 374086 105544 374092 105596
rect 374144 105584 374150 105596
rect 542354 105584 542360 105596
rect 374144 105556 542360 105584
rect 374144 105544 374150 105556
rect 542354 105544 542360 105556
rect 542412 105544 542418 105596
rect 300854 104116 300860 104168
rect 300912 104156 300918 104168
rect 375466 104156 375472 104168
rect 300912 104128 375472 104156
rect 300912 104116 300918 104128
rect 375466 104116 375472 104128
rect 375524 104116 375530 104168
rect 375558 104116 375564 104168
rect 375616 104156 375622 104168
rect 546494 104156 546500 104168
rect 375616 104128 546500 104156
rect 375616 104116 375622 104128
rect 546494 104116 546500 104128
rect 546552 104116 546558 104168
rect 378318 102756 378324 102808
rect 378376 102796 378382 102808
rect 553394 102796 553400 102808
rect 378376 102768 553400 102796
rect 378376 102756 378382 102768
rect 553394 102756 553400 102768
rect 553452 102756 553458 102808
rect 379514 101396 379520 101448
rect 379572 101436 379578 101448
rect 556246 101436 556252 101448
rect 379572 101408 556252 101436
rect 379572 101396 379578 101408
rect 556246 101396 556252 101408
rect 556304 101396 556310 101448
rect 394326 100648 394332 100700
rect 394384 100688 394390 100700
rect 580166 100688 580172 100700
rect 394384 100660 580172 100688
rect 394384 100648 394390 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 386414 98608 386420 98660
rect 386472 98648 386478 98660
rect 570598 98648 570604 98660
rect 386472 98620 570604 98648
rect 386472 98608 386478 98620
rect 570598 98608 570604 98620
rect 570656 98608 570662 98660
rect 389266 97248 389272 97300
rect 389324 97288 389330 97300
rect 578234 97288 578240 97300
rect 389324 97260 578240 97288
rect 389324 97248 389330 97260
rect 578234 97248 578240 97260
rect 578292 97248 578298 97300
rect 334066 94460 334072 94512
rect 334124 94500 334130 94512
rect 451274 94500 451280 94512
rect 334124 94472 451280 94500
rect 334124 94460 334130 94472
rect 451274 94460 451280 94472
rect 451332 94460 451338 94512
rect 327166 93100 327172 93152
rect 327224 93140 327230 93152
rect 437474 93140 437480 93152
rect 327224 93112 437480 93140
rect 327224 93100 327230 93112
rect 437474 93100 437480 93112
rect 437532 93100 437538 93152
rect 292758 91740 292764 91792
rect 292816 91780 292822 91792
rect 357526 91780 357532 91792
rect 292816 91752 357532 91780
rect 292816 91740 292822 91752
rect 357526 91740 357532 91752
rect 357584 91740 357590 91792
rect 357618 91740 357624 91792
rect 357676 91780 357682 91792
rect 505094 91780 505100 91792
rect 357676 91752 505100 91780
rect 357676 91740 357682 91752
rect 505094 91740 505100 91752
rect 505152 91740 505158 91792
rect 396718 86912 396724 86964
rect 396776 86952 396782 86964
rect 580166 86952 580172 86964
rect 396776 86924 580172 86952
rect 396776 86912 396782 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 189902 85524 189908 85536
rect 3384 85496 189908 85524
rect 3384 85484 3390 85496
rect 189902 85484 189908 85496
rect 189960 85484 189966 85536
rect 394234 73108 394240 73160
rect 394292 73148 394298 73160
rect 580166 73148 580172 73160
rect 394292 73120 580172 73148
rect 394292 73108 394298 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 21358 71720 21364 71732
rect 3384 71692 21364 71720
rect 3384 71680 3390 71692
rect 21358 71680 21364 71692
rect 21416 71680 21422 71732
rect 309134 61344 309140 61396
rect 309192 61384 309198 61396
rect 393314 61384 393320 61396
rect 309192 61356 393320 61384
rect 309192 61344 309198 61356
rect 393314 61344 393320 61356
rect 393372 61344 393378 61396
rect 394142 60664 394148 60716
rect 394200 60704 394206 60716
rect 580166 60704 580172 60716
rect 394200 60676 580172 60704
rect 394200 60664 394206 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 303706 59984 303712 60036
rect 303764 60024 303770 60036
rect 382366 60024 382372 60036
rect 303764 59996 382372 60024
rect 303764 59984 303770 59996
rect 382366 59984 382372 59996
rect 382424 59984 382430 60036
rect 305178 58624 305184 58676
rect 305236 58664 305242 58676
rect 386414 58664 386420 58676
rect 305236 58636 386420 58664
rect 305236 58624 305242 58636
rect 386414 58624 386420 58636
rect 386472 58624 386478 58676
rect 302418 57196 302424 57248
rect 302476 57236 302482 57248
rect 379514 57236 379520 57248
rect 302476 57208 379520 57236
rect 302476 57196 302482 57208
rect 379514 57196 379520 57208
rect 379572 57196 379578 57248
rect 299566 55836 299572 55888
rect 299624 55876 299630 55888
rect 372614 55876 372620 55888
rect 299624 55848 372620 55876
rect 299624 55836 299630 55848
rect 372614 55836 372620 55848
rect 372672 55836 372678 55888
rect 291378 54476 291384 54528
rect 291436 54516 291442 54528
rect 354674 54516 354680 54528
rect 291436 54488 354680 54516
rect 291436 54476 291442 54488
rect 354674 54476 354680 54488
rect 354732 54476 354738 54528
rect 296714 53048 296720 53100
rect 296772 53088 296778 53100
rect 365806 53088 365812 53100
rect 296772 53060 365812 53088
rect 296772 53048 296778 53060
rect 365806 53048 365812 53060
rect 365864 53048 365870 53100
rect 294138 51688 294144 51740
rect 294196 51728 294202 51740
rect 361574 51728 361580 51740
rect 294196 51700 361580 51728
rect 294196 51688 294202 51700
rect 361574 51688 361580 51700
rect 361632 51688 361638 51740
rect 383654 51688 383660 51740
rect 383712 51728 383718 51740
rect 566458 51728 566464 51740
rect 383712 51700 566464 51728
rect 383712 51688 383718 51700
rect 566458 51688 566464 51700
rect 566516 51688 566522 51740
rect 289814 50328 289820 50380
rect 289872 50368 289878 50380
rect 350534 50368 350540 50380
rect 289872 50340 350540 50368
rect 289872 50328 289878 50340
rect 350534 50328 350540 50340
rect 350592 50328 350598 50380
rect 295978 48968 295984 49020
rect 296036 49008 296042 49020
rect 352098 49008 352104 49020
rect 296036 48980 352104 49008
rect 296036 48968 296042 48980
rect 352098 48968 352104 48980
rect 352156 48968 352162 49020
rect 387886 48968 387892 49020
rect 387944 49008 387950 49020
rect 574094 49008 574100 49020
rect 387944 48980 574100 49008
rect 387944 48968 387950 48980
rect 574094 48968 574100 48980
rect 574152 48968 574158 49020
rect 292574 47676 292580 47728
rect 292632 47716 292638 47728
rect 357618 47716 357624 47728
rect 292632 47688 357624 47716
rect 292632 47676 292638 47688
rect 357618 47676 357624 47688
rect 357676 47676 357682 47728
rect 357434 47540 357440 47592
rect 357492 47580 357498 47592
rect 506566 47580 506572 47592
rect 357492 47552 506572 47580
rect 357492 47540 357498 47552
rect 506566 47540 506572 47552
rect 506624 47540 506630 47592
rect 457438 46860 457444 46912
rect 457496 46900 457502 46912
rect 580166 46900 580172 46912
rect 457496 46872 580172 46900
rect 457496 46860 457502 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 278866 46180 278872 46232
rect 278924 46220 278930 46232
rect 325694 46220 325700 46232
rect 278924 46192 325700 46220
rect 278924 46180 278930 46192
rect 325694 46180 325700 46192
rect 325752 46180 325758 46232
rect 335538 46180 335544 46232
rect 335596 46220 335602 46232
rect 456886 46220 456892 46232
rect 335596 46192 456892 46220
rect 335596 46180 335602 46192
rect 456886 46180 456892 46192
rect 456944 46180 456950 46232
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 189810 45540 189816 45552
rect 3568 45512 189816 45540
rect 3568 45500 3574 45512
rect 189810 45500 189816 45512
rect 189868 45500 189874 45552
rect 309870 44820 309876 44872
rect 309928 44860 309934 44872
rect 374086 44860 374092 44872
rect 309928 44832 374092 44860
rect 309928 44820 309934 44832
rect 374086 44820 374092 44832
rect 374144 44820 374150 44872
rect 380894 44820 380900 44872
rect 380952 44860 380958 44872
rect 560294 44860 560300 44872
rect 380952 44832 560300 44860
rect 380952 44820 380958 44832
rect 560294 44820 560300 44832
rect 560352 44820 560358 44872
rect 320818 43392 320824 43444
rect 320876 43432 320882 43444
rect 408494 43432 408500 43444
rect 320876 43404 408500 43432
rect 320876 43392 320882 43404
rect 408494 43392 408500 43404
rect 408552 43392 408558 43444
rect 303614 42168 303620 42220
rect 303672 42208 303678 42220
rect 382550 42208 382556 42220
rect 303672 42180 382556 42208
rect 303672 42168 303678 42180
rect 382550 42168 382556 42180
rect 382608 42168 382614 42220
rect 382458 42032 382464 42084
rect 382516 42072 382522 42084
rect 564526 42072 564532 42084
rect 382516 42044 564532 42072
rect 382516 42032 382522 42044
rect 564526 42032 564532 42044
rect 564584 42032 564590 42084
rect 277486 40672 277492 40724
rect 277544 40712 277550 40724
rect 323118 40712 323124 40724
rect 277544 40684 323124 40712
rect 277544 40672 277550 40684
rect 323118 40672 323124 40684
rect 323176 40672 323182 40724
rect 371878 40672 371884 40724
rect 371936 40712 371942 40724
rect 531314 40712 531320 40724
rect 371936 40684 531320 40712
rect 371936 40672 371942 40684
rect 531314 40672 531320 40684
rect 531372 40672 531378 40724
rect 276290 39312 276296 39364
rect 276348 39352 276354 39364
rect 318794 39352 318800 39364
rect 276348 39324 318800 39352
rect 276348 39312 276354 39324
rect 318794 39312 318800 39324
rect 318852 39312 318858 39364
rect 365714 39312 365720 39364
rect 365772 39352 365778 39364
rect 523034 39352 523040 39364
rect 365772 39324 523040 39352
rect 365772 39312 365778 39324
rect 523034 39312 523040 39324
rect 523092 39312 523098 39364
rect 273346 37884 273352 37936
rect 273404 37924 273410 37936
rect 311986 37924 311992 37936
rect 273404 37896 311992 37924
rect 273404 37884 273410 37896
rect 311986 37884 311992 37896
rect 312044 37884 312050 37936
rect 358814 37884 358820 37936
rect 358872 37924 358878 37936
rect 509234 37924 509240 37936
rect 358872 37896 509240 37924
rect 358872 37884 358878 37896
rect 509234 37884 509240 37896
rect 509292 37884 509298 37936
rect 300118 36524 300124 36576
rect 300176 36564 300182 36576
rect 349338 36564 349344 36576
rect 300176 36536 349344 36564
rect 300176 36524 300182 36536
rect 349338 36524 349344 36536
rect 349396 36524 349402 36576
rect 351914 36524 351920 36576
rect 351972 36564 351978 36576
rect 491294 36564 491300 36576
rect 351972 36536 491300 36564
rect 351972 36524 351978 36536
rect 491294 36524 491300 36536
rect 491352 36524 491358 36576
rect 271874 35164 271880 35216
rect 271932 35204 271938 35216
rect 307754 35204 307760 35216
rect 271932 35176 307760 35204
rect 271932 35164 271938 35176
rect 307754 35164 307760 35176
rect 307812 35164 307818 35216
rect 323026 35164 323032 35216
rect 323084 35204 323090 35216
rect 426434 35204 426440 35216
rect 323084 35176 426440 35204
rect 323084 35164 323090 35176
rect 426434 35164 426440 35176
rect 426492 35164 426498 35216
rect 287698 33736 287704 33788
rect 287756 33776 287762 33788
rect 335446 33776 335452 33788
rect 287756 33748 335452 33776
rect 287756 33736 287762 33748
rect 335446 33736 335452 33748
rect 335504 33736 335510 33788
rect 347038 33736 347044 33788
rect 347096 33776 347102 33788
rect 473446 33776 473452 33788
rect 347096 33748 473452 33776
rect 347096 33736 347102 33748
rect 473446 33736 473452 33748
rect 473504 33736 473510 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 190086 33096 190092 33108
rect 2924 33068 190092 33096
rect 2924 33056 2930 33068
rect 190086 33056 190092 33068
rect 190144 33056 190150 33108
rect 394050 33056 394056 33108
rect 394108 33096 394114 33108
rect 579890 33096 579896 33108
rect 394108 33068 579896 33096
rect 394108 33056 394114 33068
rect 579890 33056 579896 33068
rect 579948 33056 579954 33108
rect 278038 32444 278044 32496
rect 278096 32484 278102 32496
rect 310698 32484 310704 32496
rect 278096 32456 310704 32484
rect 278096 32444 278102 32456
rect 310698 32444 310704 32456
rect 310756 32444 310762 32496
rect 298278 32376 298284 32428
rect 298336 32416 298342 32428
rect 368474 32416 368480 32428
rect 298336 32388 368480 32416
rect 298336 32376 298342 32388
rect 368474 32376 368480 32388
rect 368532 32376 368538 32428
rect 270494 31016 270500 31068
rect 270552 31056 270558 31068
rect 305086 31056 305092 31068
rect 270552 31028 305092 31056
rect 270552 31016 270558 31028
rect 305086 31016 305092 31028
rect 305144 31016 305150 31068
rect 329190 31016 329196 31068
rect 329248 31056 329254 31068
rect 433334 31056 433340 31068
rect 329248 31028 433340 31056
rect 329248 31016 329254 31028
rect 433334 31016 433340 31028
rect 433392 31016 433398 31068
rect 254118 29588 254124 29640
rect 254176 29628 254182 29640
rect 267918 29628 267924 29640
rect 254176 29600 267924 29628
rect 254176 29588 254182 29600
rect 267918 29588 267924 29600
rect 267976 29588 267982 29640
rect 268010 29588 268016 29640
rect 268068 29628 268074 29640
rect 299566 29628 299572 29640
rect 268068 29600 299572 29628
rect 268068 29588 268074 29600
rect 299566 29588 299572 29600
rect 299624 29588 299630 29640
rect 323578 29588 323584 29640
rect 323636 29628 323642 29640
rect 415486 29628 415492 29640
rect 323636 29600 415492 29628
rect 323636 29588 323642 29600
rect 415486 29588 415492 29600
rect 415544 29588 415550 29640
rect 282270 28228 282276 28280
rect 282328 28268 282334 28280
rect 324498 28268 324504 28280
rect 282328 28240 324504 28268
rect 282328 28228 282334 28240
rect 324498 28228 324504 28240
rect 324556 28228 324562 28280
rect 331214 28228 331220 28280
rect 331272 28268 331278 28280
rect 444374 28268 444380 28280
rect 331272 28240 444380 28268
rect 331272 28228 331278 28240
rect 444374 28228 444380 28240
rect 444432 28228 444438 28280
rect 306374 26936 306380 26988
rect 306432 26976 306438 26988
rect 387886 26976 387892 26988
rect 306432 26948 387892 26976
rect 306432 26936 306438 26948
rect 387886 26936 387892 26948
rect 387944 26936 387950 26988
rect 267826 26868 267832 26920
rect 267884 26908 267890 26920
rect 300854 26908 300860 26920
rect 267884 26880 300860 26908
rect 267884 26868 267890 26880
rect 300854 26868 300860 26880
rect 300912 26868 300918 26920
rect 376754 26868 376760 26920
rect 376812 26908 376818 26920
rect 549254 26908 549260 26920
rect 376812 26880 549260 26908
rect 376812 26868 376818 26880
rect 549254 26868 549260 26880
rect 549312 26868 549318 26920
rect 266538 25508 266544 25560
rect 266596 25548 266602 25560
rect 298278 25548 298284 25560
rect 266596 25520 298284 25548
rect 266596 25508 266602 25520
rect 298278 25508 298284 25520
rect 298336 25508 298342 25560
rect 304994 25508 305000 25560
rect 305052 25548 305058 25560
rect 383654 25548 383660 25560
rect 305052 25520 383660 25548
rect 305052 25508 305058 25520
rect 383654 25508 383660 25520
rect 383712 25508 383718 25560
rect 385034 25508 385040 25560
rect 385092 25548 385098 25560
rect 569954 25548 569960 25560
rect 385092 25520 569960 25548
rect 385092 25508 385098 25520
rect 569954 25508 569960 25520
rect 570012 25508 570018 25560
rect 264974 24080 264980 24132
rect 265032 24120 265038 24132
rect 294138 24120 294144 24132
rect 265032 24092 294144 24120
rect 265032 24080 265038 24092
rect 294138 24080 294144 24092
rect 294196 24080 294202 24132
rect 302326 24080 302332 24132
rect 302384 24120 302390 24132
rect 380894 24120 380900 24132
rect 302384 24092 380900 24120
rect 302384 24080 302390 24092
rect 380894 24080 380900 24092
rect 380952 24080 380958 24132
rect 382274 24080 382280 24132
rect 382332 24120 382338 24132
rect 563054 24120 563060 24132
rect 382332 24092 563060 24120
rect 382332 24080 382338 24092
rect 563054 24080 563060 24092
rect 563112 24080 563118 24132
rect 298186 22788 298192 22840
rect 298244 22828 298250 22840
rect 370038 22828 370044 22840
rect 298244 22800 370044 22828
rect 298244 22788 298250 22800
rect 370038 22788 370044 22800
rect 370096 22788 370102 22840
rect 267734 22720 267740 22772
rect 267792 22760 267798 22772
rect 299658 22760 299664 22772
rect 267792 22732 299664 22760
rect 267792 22720 267798 22732
rect 299658 22720 299664 22732
rect 299716 22720 299722 22772
rect 359458 22720 359464 22772
rect 359516 22760 359522 22772
rect 498194 22760 498200 22772
rect 359516 22732 498200 22760
rect 359516 22720 359522 22732
rect 498194 22720 498200 22732
rect 498252 22720 498258 22772
rect 270678 21428 270684 21480
rect 270736 21468 270742 21480
rect 307846 21468 307852 21480
rect 270736 21440 307852 21468
rect 270736 21428 270742 21440
rect 307846 21428 307852 21440
rect 307904 21428 307910 21480
rect 284386 21360 284392 21412
rect 284444 21400 284450 21412
rect 336826 21400 336832 21412
rect 284444 21372 336832 21400
rect 284444 21360 284450 21372
rect 336826 21360 336832 21372
rect 336884 21360 336890 21412
rect 353386 21360 353392 21412
rect 353444 21400 353450 21412
rect 498286 21400 498292 21412
rect 353444 21372 498292 21400
rect 353444 21360 353450 21372
rect 498286 21360 498292 21372
rect 498344 21360 498350 21412
rect 393958 20612 393964 20664
rect 394016 20652 394022 20664
rect 579890 20652 579896 20664
rect 394016 20624 579896 20652
rect 394016 20612 394022 20624
rect 579890 20612 579896 20624
rect 579948 20612 579954 20664
rect 280246 20000 280252 20052
rect 280304 20040 280310 20052
rect 327166 20040 327172 20052
rect 280304 20012 327172 20040
rect 280304 20000 280310 20012
rect 327166 20000 327172 20012
rect 327224 20000 327230 20052
rect 310606 19932 310612 19984
rect 310664 19972 310670 19984
rect 397454 19972 397460 19984
rect 310664 19944 397460 19972
rect 310664 19932 310670 19944
rect 397454 19932 397460 19944
rect 397512 19932 397518 19984
rect 256786 18776 256792 18828
rect 256844 18816 256850 18828
rect 276198 18816 276204 18828
rect 256844 18788 276204 18816
rect 256844 18776 256850 18788
rect 276198 18776 276204 18788
rect 276256 18776 276262 18828
rect 276106 18640 276112 18692
rect 276164 18680 276170 18692
rect 320358 18680 320364 18692
rect 276164 18652 320364 18680
rect 276164 18640 276170 18652
rect 320358 18640 320364 18652
rect 320416 18640 320422 18692
rect 338758 18640 338764 18692
rect 338816 18680 338822 18692
rect 390646 18680 390652 18692
rect 338816 18652 390652 18680
rect 338816 18640 338822 18652
rect 390646 18640 390652 18652
rect 390704 18640 390710 18692
rect 287146 18572 287152 18624
rect 287204 18612 287210 18624
rect 343726 18612 343732 18624
rect 287204 18584 343732 18612
rect 287204 18572 287210 18584
rect 343726 18572 343732 18584
rect 343784 18572 343790 18624
rect 368566 18572 368572 18624
rect 368624 18612 368630 18624
rect 531406 18612 531412 18624
rect 368624 18584 531412 18612
rect 368624 18572 368630 18584
rect 531406 18572 531412 18584
rect 531464 18572 531470 18624
rect 304258 17280 304264 17332
rect 304316 17320 304322 17332
rect 365714 17320 365720 17332
rect 304316 17292 365720 17320
rect 304316 17280 304322 17292
rect 365714 17280 365720 17292
rect 365772 17280 365778 17332
rect 266354 17212 266360 17264
rect 266412 17252 266418 17264
rect 295518 17252 295524 17264
rect 266412 17224 295524 17252
rect 266412 17212 266418 17224
rect 295518 17212 295524 17224
rect 295576 17212 295582 17264
rect 364518 17212 364524 17264
rect 364576 17252 364582 17264
rect 523126 17252 523132 17264
rect 364576 17224 523132 17252
rect 364576 17212 364582 17224
rect 523126 17212 523132 17224
rect 523184 17212 523190 17264
rect 273898 15920 273904 15972
rect 273956 15960 273962 15972
rect 309686 15960 309692 15972
rect 273956 15932 309692 15960
rect 273956 15920 273962 15932
rect 309686 15920 309692 15932
rect 309744 15920 309750 15972
rect 282914 15852 282920 15904
rect 282972 15892 282978 15904
rect 332686 15892 332692 15904
rect 282972 15864 332692 15892
rect 282972 15852 282978 15864
rect 332686 15852 332692 15864
rect 332744 15852 332750 15904
rect 349430 15852 349436 15904
rect 349488 15892 349494 15904
rect 487154 15892 487160 15904
rect 349488 15864 487160 15892
rect 349488 15852 349494 15864
rect 487154 15852 487160 15864
rect 487212 15852 487218 15904
rect 270586 14492 270592 14544
rect 270644 14532 270650 14544
rect 306374 14532 306380 14544
rect 270644 14504 306380 14532
rect 270644 14492 270650 14504
rect 306374 14492 306380 14504
rect 306432 14492 306438 14544
rect 309778 14492 309784 14544
rect 309836 14532 309842 14544
rect 390922 14532 390928 14544
rect 309836 14504 390928 14532
rect 309836 14492 309842 14504
rect 390922 14492 390928 14504
rect 390980 14492 390986 14544
rect 274726 14424 274732 14476
rect 274784 14464 274790 14476
rect 316218 14464 316224 14476
rect 274784 14436 316224 14464
rect 274784 14424 274790 14436
rect 316218 14424 316224 14436
rect 316276 14424 316282 14476
rect 346486 14424 346492 14476
rect 346544 14464 346550 14476
rect 480530 14464 480536 14476
rect 346544 14436 480536 14464
rect 346544 14424 346550 14436
rect 480530 14424 480536 14436
rect 480588 14424 480594 14476
rect 356146 13268 356152 13320
rect 356204 13308 356210 13320
rect 503714 13308 503720 13320
rect 356204 13280 503720 13308
rect 356204 13268 356210 13280
rect 503714 13268 503720 13280
rect 503772 13268 503778 13320
rect 340966 13200 340972 13252
rect 341024 13240 341030 13252
rect 341150 13240 341156 13252
rect 341024 13212 341156 13240
rect 341024 13200 341030 13212
rect 341150 13200 341156 13212
rect 341208 13200 341214 13252
rect 360194 13200 360200 13252
rect 360252 13240 360258 13252
rect 511258 13240 511264 13252
rect 360252 13212 511264 13240
rect 360252 13200 360258 13212
rect 511258 13200 511264 13212
rect 511316 13200 511322 13252
rect 266446 13132 266452 13184
rect 266504 13172 266510 13184
rect 297266 13172 297272 13184
rect 266504 13144 297272 13172
rect 266504 13132 266510 13144
rect 297266 13132 297272 13144
rect 297324 13132 297330 13184
rect 363046 13132 363052 13184
rect 363104 13172 363110 13184
rect 517882 13172 517888 13184
rect 363104 13144 517888 13172
rect 363104 13132 363110 13144
rect 517882 13132 517888 13144
rect 517940 13132 517946 13184
rect 197906 13064 197912 13116
rect 197964 13104 197970 13116
rect 222286 13104 222292 13116
rect 197964 13076 222292 13104
rect 197964 13064 197970 13076
rect 222286 13064 222292 13076
rect 222344 13064 222350 13116
rect 254026 13064 254032 13116
rect 254084 13104 254090 13116
rect 267734 13104 267740 13116
rect 254084 13076 267740 13104
rect 254084 13064 254090 13076
rect 267734 13064 267740 13076
rect 267792 13064 267798 13116
rect 269206 13064 269212 13116
rect 269264 13104 269270 13116
rect 303154 13104 303160 13116
rect 269264 13076 303160 13104
rect 269264 13064 269270 13076
rect 303154 13064 303160 13076
rect 303212 13064 303218 13116
rect 307018 13064 307024 13116
rect 307076 13104 307082 13116
rect 340966 13104 340972 13116
rect 307076 13076 340972 13104
rect 307076 13064 307082 13076
rect 340966 13064 340972 13076
rect 341024 13064 341030 13116
rect 364426 13064 364432 13116
rect 364484 13104 364490 13116
rect 521654 13104 521660 13116
rect 364484 13076 521660 13104
rect 364484 13064 364490 13076
rect 521654 13064 521660 13076
rect 521712 13064 521718 13116
rect 341058 12044 341064 12096
rect 341116 12084 341122 12096
rect 467466 12084 467472 12096
rect 341116 12056 467472 12084
rect 341116 12044 341122 12056
rect 467466 12044 467472 12056
rect 467524 12044 467530 12096
rect 342346 11976 342352 12028
rect 342404 12016 342410 12028
rect 470594 12016 470600 12028
rect 342404 11988 470600 12016
rect 342404 11976 342410 11988
rect 470594 11976 470600 11988
rect 470652 11976 470658 12028
rect 345198 11908 345204 11960
rect 345256 11948 345262 11960
rect 478138 11948 478144 11960
rect 345256 11920 478144 11948
rect 345256 11908 345262 11920
rect 478138 11908 478144 11920
rect 478196 11908 478202 11960
rect 259638 11840 259644 11892
rect 259696 11880 259702 11892
rect 281626 11880 281632 11892
rect 259696 11852 281632 11880
rect 259696 11840 259702 11852
rect 281626 11840 281632 11852
rect 281684 11840 281690 11892
rect 349246 11840 349252 11892
rect 349304 11880 349310 11892
rect 486418 11880 486424 11892
rect 349304 11852 486424 11880
rect 349304 11840 349310 11852
rect 486418 11840 486424 11852
rect 486476 11840 486482 11892
rect 176654 11772 176660 11824
rect 176712 11812 176718 11824
rect 177850 11812 177856 11824
rect 176712 11784 177856 11812
rect 176712 11772 176718 11784
rect 177850 11772 177856 11784
rect 177908 11772 177914 11824
rect 201494 11772 201500 11824
rect 201552 11812 201558 11824
rect 202690 11812 202696 11824
rect 201552 11784 202696 11812
rect 201552 11772 201558 11784
rect 202690 11772 202696 11784
rect 202748 11772 202754 11824
rect 273254 11772 273260 11824
rect 273312 11812 273318 11824
rect 313826 11812 313832 11824
rect 273312 11784 313832 11812
rect 273312 11772 273318 11784
rect 313826 11772 313832 11784
rect 313884 11772 313890 11824
rect 352006 11772 352012 11824
rect 352064 11812 352070 11824
rect 493042 11812 493048 11824
rect 352064 11784 493048 11812
rect 352064 11772 352070 11784
rect 493042 11772 493048 11784
rect 493100 11772 493106 11824
rect 169570 11704 169576 11756
rect 169628 11744 169634 11756
rect 209866 11744 209872 11756
rect 169628 11716 209872 11744
rect 169628 11704 169634 11716
rect 209866 11704 209872 11716
rect 209924 11704 209930 11756
rect 242894 11704 242900 11756
rect 242952 11744 242958 11756
rect 244090 11744 244096 11756
rect 242952 11716 244096 11744
rect 242952 11704 242958 11716
rect 244090 11704 244096 11716
rect 244148 11704 244154 11756
rect 281534 11704 281540 11756
rect 281592 11744 281598 11756
rect 281592 11716 316034 11744
rect 281592 11704 281598 11716
rect 316006 11676 316034 11716
rect 329098 11704 329104 11756
rect 329156 11744 329162 11756
rect 331214 11744 331220 11756
rect 329156 11716 331220 11744
rect 329156 11704 329162 11716
rect 331214 11704 331220 11716
rect 331272 11704 331278 11756
rect 353294 11704 353300 11756
rect 353352 11744 353358 11756
rect 497090 11744 497096 11756
rect 353352 11716 497096 11744
rect 353352 11704 353358 11716
rect 497090 11704 497096 11716
rect 497148 11704 497154 11756
rect 332778 11676 332784 11688
rect 316006 11648 332784 11676
rect 332778 11636 332784 11648
rect 332836 11636 332842 11688
rect 310514 10684 310520 10736
rect 310572 10724 310578 10736
rect 398926 10724 398932 10736
rect 310572 10696 398932 10724
rect 310572 10684 310578 10696
rect 398926 10684 398932 10696
rect 398984 10684 398990 10736
rect 313274 10616 313280 10668
rect 313332 10656 313338 10668
rect 403618 10656 403624 10668
rect 313332 10628 403624 10656
rect 313332 10616 313338 10628
rect 403618 10616 403624 10628
rect 403676 10616 403682 10668
rect 316126 10548 316132 10600
rect 316184 10588 316190 10600
rect 410794 10588 410800 10600
rect 316184 10560 410800 10588
rect 316184 10548 316190 10560
rect 410794 10548 410800 10560
rect 410852 10548 410858 10600
rect 201678 10480 201684 10532
rect 201736 10520 201742 10532
rect 209038 10520 209044 10532
rect 201736 10492 209044 10520
rect 201736 10480 201742 10492
rect 209038 10480 209044 10492
rect 209096 10480 209102 10532
rect 317598 10480 317604 10532
rect 317656 10520 317662 10532
rect 414290 10520 414296 10532
rect 317656 10492 414296 10520
rect 317656 10480 317662 10492
rect 414290 10480 414296 10492
rect 414348 10480 414354 10532
rect 262490 10412 262496 10464
rect 262548 10452 262554 10464
rect 288986 10452 288992 10464
rect 262548 10424 288992 10452
rect 262548 10412 262554 10424
rect 288986 10412 288992 10424
rect 289044 10412 289050 10464
rect 320266 10412 320272 10464
rect 320324 10452 320330 10464
rect 420914 10452 420920 10464
rect 320324 10424 420920 10452
rect 320324 10412 320330 10424
rect 420914 10412 420920 10424
rect 420972 10412 420978 10464
rect 263778 10344 263784 10396
rect 263836 10384 263842 10396
rect 289814 10384 289820 10396
rect 263836 10356 289820 10384
rect 263836 10344 263842 10356
rect 289814 10344 289820 10356
rect 289872 10344 289878 10396
rect 321646 10344 321652 10396
rect 321704 10384 321710 10396
rect 423766 10384 423772 10396
rect 321704 10356 423772 10384
rect 321704 10344 321710 10356
rect 423766 10344 423772 10356
rect 423824 10344 423830 10396
rect 128998 10276 129004 10328
rect 129056 10316 129062 10328
rect 191926 10316 191932 10328
rect 129056 10288 191932 10316
rect 129056 10276 129062 10288
rect 191926 10276 191932 10288
rect 191984 10276 191990 10328
rect 207106 10276 207112 10328
rect 207164 10316 207170 10328
rect 226978 10316 226984 10328
rect 207164 10288 226984 10316
rect 207164 10276 207170 10288
rect 226978 10276 226984 10288
rect 227036 10276 227042 10328
rect 274634 10276 274640 10328
rect 274692 10316 274698 10328
rect 314654 10316 314660 10328
rect 274692 10288 314660 10316
rect 274692 10276 274698 10288
rect 314654 10276 314660 10288
rect 314712 10276 314718 10328
rect 322934 10276 322940 10328
rect 322992 10316 322998 10328
rect 428458 10316 428464 10328
rect 322992 10288 428464 10316
rect 322992 10276 322998 10288
rect 428458 10276 428464 10288
rect 428516 10276 428522 10328
rect 302234 9324 302240 9376
rect 302292 9364 302298 9376
rect 378870 9364 378876 9376
rect 302292 9336 378876 9364
rect 302292 9324 302298 9336
rect 378870 9324 378876 9336
rect 378928 9324 378934 9376
rect 367094 9256 367100 9308
rect 367152 9296 367158 9308
rect 527818 9296 527824 9308
rect 367152 9268 527824 9296
rect 367152 9256 367158 9268
rect 527818 9256 527824 9268
rect 527876 9256 527882 9308
rect 369946 9188 369952 9240
rect 370004 9228 370010 9240
rect 534902 9228 534908 9240
rect 370004 9200 534908 9228
rect 370004 9188 370010 9200
rect 534902 9188 534908 9200
rect 534960 9188 534966 9240
rect 291286 9120 291292 9172
rect 291344 9160 291350 9172
rect 354030 9160 354036 9172
rect 291344 9132 354036 9160
rect 291344 9120 291350 9132
rect 354030 9120 354036 9132
rect 354088 9120 354094 9172
rect 371326 9120 371332 9172
rect 371384 9160 371390 9172
rect 538398 9160 538404 9172
rect 371384 9132 538404 9160
rect 371384 9120 371390 9132
rect 538398 9120 538404 9132
rect 538456 9120 538462 9172
rect 294046 9052 294052 9104
rect 294104 9092 294110 9104
rect 361114 9092 361120 9104
rect 294104 9064 361120 9092
rect 294104 9052 294110 9064
rect 361114 9052 361120 9064
rect 361172 9052 361178 9104
rect 373994 9052 374000 9104
rect 374052 9092 374058 9104
rect 545482 9092 545488 9104
rect 374052 9064 545488 9092
rect 374052 9052 374058 9064
rect 545482 9052 545488 9064
rect 545540 9052 545546 9104
rect 258350 8984 258356 9036
rect 258408 9024 258414 9036
rect 278314 9024 278320 9036
rect 258408 8996 278320 9024
rect 258408 8984 258414 8996
rect 278314 8984 278320 8996
rect 278372 8984 278378 9036
rect 282178 8984 282184 9036
rect 282236 9024 282242 9036
rect 293678 9024 293684 9036
rect 282236 8996 293684 9024
rect 282236 8984 282242 8996
rect 293678 8984 293684 8996
rect 293736 8984 293742 9036
rect 295426 8984 295432 9036
rect 295484 9024 295490 9036
rect 364610 9024 364616 9036
rect 295484 8996 364616 9024
rect 295484 8984 295490 8996
rect 364610 8984 364616 8996
rect 364668 8984 364674 9036
rect 375374 8984 375380 9036
rect 375432 9024 375438 9036
rect 549070 9024 549076 9036
rect 375432 8996 549076 9024
rect 375432 8984 375438 8996
rect 549070 8984 549076 8996
rect 549128 8984 549134 9036
rect 154206 8916 154212 8968
rect 154264 8956 154270 8968
rect 188338 8956 188344 8968
rect 154264 8928 188344 8956
rect 154264 8916 154270 8928
rect 188338 8916 188344 8928
rect 188396 8916 188402 8968
rect 200298 8916 200304 8968
rect 200356 8956 200362 8968
rect 223666 8956 223672 8968
rect 200356 8928 223672 8956
rect 200356 8916 200362 8928
rect 223666 8916 223672 8928
rect 223724 8916 223730 8968
rect 263686 8916 263692 8968
rect 263744 8956 263750 8968
rect 292574 8956 292580 8968
rect 263744 8928 292580 8956
rect 263744 8916 263750 8928
rect 292574 8916 292580 8928
rect 292632 8916 292638 8968
rect 298094 8916 298100 8968
rect 298152 8956 298158 8968
rect 371694 8956 371700 8968
rect 298152 8928 371700 8956
rect 298152 8916 298158 8928
rect 371694 8916 371700 8928
rect 371752 8916 371758 8968
rect 378134 8916 378140 8968
rect 378192 8956 378198 8968
rect 552658 8956 552664 8968
rect 378192 8928 552664 8956
rect 378192 8916 378198 8928
rect 552658 8916 552664 8928
rect 552716 8916 552722 8968
rect 288526 8032 288532 8084
rect 288584 8072 288590 8084
rect 346946 8072 346952 8084
rect 288584 8044 346952 8072
rect 288584 8032 288590 8044
rect 346946 8032 346952 8044
rect 347004 8032 347010 8084
rect 335354 7964 335360 8016
rect 335412 8004 335418 8016
rect 455690 8004 455696 8016
rect 335412 7976 455696 8004
rect 335412 7964 335418 7976
rect 455690 7964 455696 7976
rect 455748 7964 455754 8016
rect 338114 7896 338120 7948
rect 338172 7936 338178 7948
rect 462774 7936 462780 7948
rect 338172 7908 462780 7936
rect 338172 7896 338178 7908
rect 462774 7896 462780 7908
rect 462832 7896 462838 7948
rect 339678 7828 339684 7880
rect 339736 7868 339742 7880
rect 466270 7868 466276 7880
rect 339736 7840 466276 7868
rect 339736 7828 339742 7840
rect 466270 7828 466276 7840
rect 466328 7828 466334 7880
rect 341150 7760 341156 7812
rect 341208 7800 341214 7812
rect 469858 7800 469864 7812
rect 341208 7772 469864 7800
rect 341208 7760 341214 7772
rect 469858 7760 469864 7772
rect 469916 7760 469922 7812
rect 345106 7692 345112 7744
rect 345164 7732 345170 7744
rect 476942 7732 476948 7744
rect 345164 7704 476948 7732
rect 345164 7692 345170 7704
rect 476942 7692 476948 7704
rect 477000 7692 477006 7744
rect 194410 7624 194416 7676
rect 194468 7664 194474 7676
rect 217318 7664 217324 7676
rect 194468 7636 217324 7664
rect 194468 7624 194474 7636
rect 217318 7624 217324 7636
rect 217376 7624 217382 7676
rect 256694 7624 256700 7676
rect 256752 7664 256758 7676
rect 274818 7664 274824 7676
rect 256752 7636 274824 7664
rect 256752 7624 256758 7636
rect 274818 7624 274824 7636
rect 274876 7624 274882 7676
rect 284478 7624 284484 7676
rect 284536 7664 284542 7676
rect 339862 7664 339868 7676
rect 284536 7636 339868 7664
rect 284536 7624 284542 7636
rect 339862 7624 339868 7636
rect 339920 7624 339926 7676
rect 346394 7624 346400 7676
rect 346452 7664 346458 7676
rect 481726 7664 481732 7676
rect 346452 7636 481732 7664
rect 346452 7624 346458 7636
rect 481726 7624 481732 7636
rect 481784 7624 481790 7676
rect 171962 7556 171968 7608
rect 172020 7596 172026 7608
rect 191098 7596 191104 7608
rect 172020 7568 191104 7596
rect 172020 7556 172026 7568
rect 191098 7556 191104 7568
rect 191156 7556 191162 7608
rect 196802 7556 196808 7608
rect 196860 7596 196866 7608
rect 222194 7596 222200 7608
rect 196860 7568 222200 7596
rect 196860 7556 196866 7568
rect 222194 7556 222200 7568
rect 222252 7556 222258 7608
rect 259546 7556 259552 7608
rect 259604 7596 259610 7608
rect 283098 7596 283104 7608
rect 259604 7568 283104 7596
rect 259604 7556 259610 7568
rect 283098 7556 283104 7568
rect 283156 7556 283162 7608
rect 285858 7556 285864 7608
rect 285916 7596 285922 7608
rect 343358 7596 343364 7608
rect 285916 7568 343364 7596
rect 285916 7556 285922 7568
rect 343358 7556 343364 7568
rect 343416 7556 343422 7608
rect 349154 7556 349160 7608
rect 349212 7596 349218 7608
rect 488810 7596 488816 7608
rect 349212 7568 488816 7596
rect 349212 7556 349218 7568
rect 488810 7556 488816 7568
rect 488868 7556 488874 7608
rect 374086 7488 374092 7540
rect 374144 7528 374150 7540
rect 375282 7528 375288 7540
rect 374144 7500 375288 7528
rect 374144 7488 374150 7500
rect 375282 7488 375288 7500
rect 375340 7488 375346 7540
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 189718 6848 189724 6860
rect 3476 6820 189724 6848
rect 3476 6808 3482 6820
rect 189718 6808 189724 6820
rect 189776 6808 189782 6860
rect 576118 6808 576124 6860
rect 576176 6848 576182 6860
rect 580166 6848 580172 6860
rect 576176 6820 580172 6848
rect 576176 6808 576182 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 276106 6536 276112 6588
rect 276164 6576 276170 6588
rect 318518 6576 318524 6588
rect 276164 6548 318524 6576
rect 276164 6536 276170 6548
rect 318518 6536 318524 6548
rect 318576 6536 318582 6588
rect 277394 6468 277400 6520
rect 277452 6508 277458 6520
rect 322106 6508 322112 6520
rect 277452 6480 322112 6508
rect 277452 6468 277458 6480
rect 322106 6468 322112 6480
rect 322164 6468 322170 6520
rect 311894 6400 311900 6452
rect 311952 6440 311958 6452
rect 402514 6440 402520 6452
rect 311952 6412 402520 6440
rect 311952 6400 311958 6412
rect 402514 6400 402520 6412
rect 402572 6400 402578 6452
rect 313366 6332 313372 6384
rect 313424 6372 313430 6384
rect 406010 6372 406016 6384
rect 313424 6344 406016 6372
rect 313424 6332 313430 6344
rect 406010 6332 406016 6344
rect 406068 6332 406074 6384
rect 203886 6264 203892 6316
rect 203944 6304 203950 6316
rect 214558 6304 214564 6316
rect 203944 6276 214564 6304
rect 203944 6264 203950 6276
rect 214558 6264 214564 6276
rect 214616 6264 214622 6316
rect 317414 6264 317420 6316
rect 317472 6304 317478 6316
rect 413094 6304 413100 6316
rect 317472 6276 413100 6304
rect 317472 6264 317478 6276
rect 413094 6264 413100 6276
rect 413152 6264 413158 6316
rect 214466 6196 214472 6248
rect 214524 6236 214530 6248
rect 230566 6236 230572 6248
rect 214524 6208 230572 6236
rect 214524 6196 214530 6208
rect 230566 6196 230572 6208
rect 230624 6196 230630 6248
rect 250070 6196 250076 6248
rect 250128 6236 250134 6248
rect 260650 6236 260656 6248
rect 250128 6208 260656 6236
rect 250128 6196 250134 6208
rect 260650 6196 260656 6208
rect 260708 6196 260714 6248
rect 269114 6196 269120 6248
rect 269172 6236 269178 6248
rect 304350 6236 304356 6248
rect 269172 6208 304356 6236
rect 269172 6196 269178 6208
rect 304350 6196 304356 6208
rect 304408 6196 304414 6248
rect 320174 6196 320180 6248
rect 320232 6236 320238 6248
rect 420178 6236 420184 6248
rect 320232 6208 420184 6236
rect 320232 6196 320238 6208
rect 420178 6196 420184 6208
rect 420236 6196 420242 6248
rect 186130 6128 186136 6180
rect 186188 6168 186194 6180
rect 216950 6168 216956 6180
rect 186188 6140 216956 6168
rect 186188 6128 186194 6140
rect 216950 6128 216956 6140
rect 217008 6128 217014 6180
rect 255498 6128 255504 6180
rect 255556 6168 255562 6180
rect 272426 6168 272432 6180
rect 255556 6140 272432 6168
rect 255556 6128 255562 6140
rect 272426 6128 272432 6140
rect 272484 6128 272490 6180
rect 280154 6128 280160 6180
rect 280212 6168 280218 6180
rect 329190 6168 329196 6180
rect 280212 6140 329196 6168
rect 280212 6128 280218 6140
rect 329190 6128 329196 6140
rect 329248 6128 329254 6180
rect 387794 6128 387800 6180
rect 387852 6168 387858 6180
rect 576302 6168 576308 6180
rect 387852 6140 576308 6168
rect 387852 6128 387858 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 189718 5244 189724 5296
rect 189776 5284 189782 5296
rect 219526 5284 219532 5296
rect 189776 5256 219532 5284
rect 189776 5244 189782 5256
rect 219526 5244 219532 5256
rect 219584 5244 219590 5296
rect 182542 5176 182548 5228
rect 182600 5216 182606 5228
rect 215570 5216 215576 5228
rect 182600 5188 215576 5216
rect 182600 5176 182606 5188
rect 215570 5176 215576 5188
rect 215628 5176 215634 5228
rect 284294 5176 284300 5228
rect 284352 5216 284358 5228
rect 338666 5216 338672 5228
rect 284352 5188 338672 5216
rect 284352 5176 284358 5188
rect 338666 5176 338672 5188
rect 338724 5176 338730 5228
rect 390738 5176 390744 5228
rect 390796 5216 390802 5228
rect 391014 5216 391020 5228
rect 390796 5188 391020 5216
rect 390796 5176 390802 5188
rect 391014 5176 391020 5188
rect 391072 5176 391078 5228
rect 179046 5108 179052 5160
rect 179104 5148 179110 5160
rect 214098 5148 214104 5160
rect 179104 5120 214104 5148
rect 179104 5108 179110 5120
rect 214098 5108 214104 5120
rect 214156 5108 214162 5160
rect 285766 5108 285772 5160
rect 285824 5148 285830 5160
rect 342162 5148 342168 5160
rect 285824 5120 342168 5148
rect 285824 5108 285830 5120
rect 342162 5108 342168 5120
rect 342220 5108 342226 5160
rect 175458 5040 175464 5092
rect 175516 5080 175522 5092
rect 212626 5080 212632 5092
rect 175516 5052 212632 5080
rect 175516 5040 175522 5052
rect 212626 5040 212632 5052
rect 212684 5040 212690 5092
rect 299474 5040 299480 5092
rect 299532 5080 299538 5092
rect 373994 5080 374000 5092
rect 299532 5052 374000 5080
rect 299532 5040 299538 5052
rect 373994 5040 374000 5052
rect 374052 5040 374058 5092
rect 140130 4972 140136 5024
rect 140188 5012 140194 5024
rect 197446 5012 197452 5024
rect 140188 4984 197452 5012
rect 140188 4972 140194 4984
rect 197446 4972 197452 4984
rect 197504 4972 197510 5024
rect 287054 4972 287060 5024
rect 287112 5012 287118 5024
rect 345750 5012 345756 5024
rect 287112 4984 345756 5012
rect 287112 4972 287118 4984
rect 345750 4972 345756 4984
rect 345808 4972 345814 5024
rect 360286 4972 360292 5024
rect 360344 5012 360350 5024
rect 512454 5012 512460 5024
rect 360344 4984 512460 5012
rect 360344 4972 360350 4984
rect 512454 4972 512460 4984
rect 512512 4972 512518 5024
rect 519538 5012 519544 5024
rect 518866 4984 519544 5012
rect 136450 4904 136456 4956
rect 136508 4944 136514 4956
rect 195974 4944 195980 4956
rect 136508 4916 195980 4944
rect 136508 4904 136514 4916
rect 195974 4904 195980 4916
rect 196032 4904 196038 4956
rect 269758 4904 269764 4956
rect 269816 4944 269822 4956
rect 285398 4944 285404 4956
rect 269816 4916 285404 4944
rect 269816 4904 269822 4916
rect 285398 4904 285404 4916
rect 285456 4904 285462 4956
rect 288434 4904 288440 4956
rect 288492 4944 288498 4956
rect 349246 4944 349252 4956
rect 288492 4916 349252 4944
rect 288492 4904 288498 4916
rect 349246 4904 349252 4916
rect 349304 4904 349310 4956
rect 362954 4904 362960 4956
rect 363012 4944 363018 4956
rect 518866 4944 518894 4984
rect 519538 4972 519544 4984
rect 519596 4972 519602 5024
rect 363012 4916 518894 4944
rect 363012 4904 363018 4916
rect 132954 4836 132960 4888
rect 133012 4876 133018 4888
rect 194778 4876 194784 4888
rect 133012 4848 194784 4876
rect 133012 4836 133018 4848
rect 194778 4836 194784 4848
rect 194836 4836 194842 4888
rect 218054 4836 218060 4888
rect 218112 4876 218118 4888
rect 232038 4876 232044 4888
rect 218112 4848 232044 4876
rect 218112 4836 218118 4848
rect 232038 4836 232044 4848
rect 232096 4836 232102 4888
rect 255406 4836 255412 4888
rect 255464 4876 255470 4888
rect 271230 4876 271236 4888
rect 255464 4848 271236 4876
rect 255464 4836 255470 4848
rect 271230 4836 271236 4848
rect 271288 4836 271294 4888
rect 293954 4836 293960 4888
rect 294012 4876 294018 4888
rect 359918 4876 359924 4888
rect 294012 4848 359924 4876
rect 294012 4836 294018 4848
rect 359918 4836 359924 4848
rect 359976 4836 359982 4888
rect 369854 4836 369860 4888
rect 369912 4876 369918 4888
rect 533706 4876 533712 4888
rect 369912 4848 533712 4876
rect 369912 4836 369918 4848
rect 533706 4836 533712 4848
rect 533764 4836 533770 4888
rect 129366 4768 129372 4820
rect 129424 4808 129430 4820
rect 193306 4808 193312 4820
rect 129424 4780 193312 4808
rect 129424 4768 129430 4780
rect 193306 4768 193312 4780
rect 193364 4768 193370 4820
rect 220906 4808 220912 4820
rect 200086 4780 220912 4808
rect 193214 4700 193220 4752
rect 193272 4740 193278 4752
rect 200086 4740 200114 4780
rect 220906 4768 220912 4780
rect 220964 4768 220970 4820
rect 258258 4768 258264 4820
rect 258316 4808 258322 4820
rect 279510 4808 279516 4820
rect 258316 4780 279516 4808
rect 258316 4768 258322 4780
rect 279510 4768 279516 4780
rect 279568 4768 279574 4820
rect 295334 4768 295340 4820
rect 295392 4808 295398 4820
rect 363506 4808 363512 4820
rect 295392 4780 363512 4808
rect 295392 4768 295398 4780
rect 363506 4768 363512 4780
rect 363564 4768 363570 4820
rect 371234 4768 371240 4820
rect 371292 4808 371298 4820
rect 537202 4808 537208 4820
rect 371292 4780 537208 4808
rect 371292 4768 371298 4780
rect 537202 4768 537208 4780
rect 537260 4768 537266 4820
rect 193272 4712 200114 4740
rect 193272 4700 193278 4712
rect 141234 4088 141240 4140
rect 141292 4128 141298 4140
rect 142798 4128 142804 4140
rect 141292 4100 142804 4128
rect 141292 4088 141298 4100
rect 142798 4088 142804 4100
rect 142856 4088 142862 4140
rect 174262 4088 174268 4140
rect 174320 4128 174326 4140
rect 212534 4128 212540 4140
rect 174320 4100 212540 4128
rect 174320 4088 174326 4100
rect 212534 4088 212540 4100
rect 212592 4088 212598 4140
rect 219250 4088 219256 4140
rect 219308 4128 219314 4140
rect 232130 4128 232136 4140
rect 219308 4100 232136 4128
rect 219308 4088 219314 4100
rect 232130 4088 232136 4100
rect 232188 4088 232194 4140
rect 251174 4088 251180 4140
rect 251232 4128 251238 4140
rect 261754 4128 261760 4140
rect 251232 4100 261760 4128
rect 251232 4088 251238 4100
rect 261754 4088 261760 4100
rect 261812 4088 261818 4140
rect 327074 4088 327080 4140
rect 327132 4128 327138 4140
rect 436738 4128 436744 4140
rect 327132 4100 436744 4128
rect 327132 4088 327138 4100
rect 436738 4088 436744 4100
rect 436796 4088 436802 4140
rect 566458 4088 566464 4140
rect 566516 4128 566522 4140
rect 568022 4128 568028 4140
rect 566516 4100 568028 4128
rect 566516 4088 566522 4100
rect 568022 4088 568028 4100
rect 568080 4088 568086 4140
rect 128170 4020 128176 4072
rect 128228 4060 128234 4072
rect 134518 4060 134524 4072
rect 128228 4032 134524 4060
rect 128228 4020 128234 4032
rect 134518 4020 134524 4032
rect 134576 4020 134582 4072
rect 167178 4020 167184 4072
rect 167236 4060 167242 4072
rect 208578 4060 208584 4072
rect 167236 4032 208584 4060
rect 167236 4020 167242 4032
rect 208578 4020 208584 4032
rect 208636 4020 208642 4072
rect 220446 4020 220452 4072
rect 220504 4060 220510 4072
rect 233234 4060 233240 4072
rect 220504 4032 233240 4060
rect 220504 4020 220510 4032
rect 233234 4020 233240 4032
rect 233292 4020 233298 4072
rect 329926 4020 329932 4072
rect 329984 4060 329990 4072
rect 443822 4060 443828 4072
rect 329984 4032 443828 4060
rect 329984 4020 329990 4032
rect 443822 4020 443828 4032
rect 443880 4020 443886 4072
rect 170766 3952 170772 4004
rect 170824 3992 170830 4004
rect 211338 3992 211344 4004
rect 170824 3964 211344 3992
rect 170824 3952 170830 3964
rect 211338 3952 211344 3964
rect 211396 3952 211402 4004
rect 215662 3952 215668 4004
rect 215720 3992 215726 4004
rect 230474 3992 230480 4004
rect 215720 3964 230480 3992
rect 215720 3952 215726 3964
rect 230474 3952 230480 3964
rect 230532 3952 230538 4004
rect 332594 3952 332600 4004
rect 332652 3992 332658 4004
rect 450906 3992 450912 4004
rect 332652 3964 450912 3992
rect 332652 3952 332658 3964
rect 450906 3952 450912 3964
rect 450964 3952 450970 4004
rect 163682 3884 163688 3936
rect 163740 3924 163746 3936
rect 207198 3924 207204 3936
rect 163740 3896 207204 3924
rect 163740 3884 163746 3896
rect 207198 3884 207204 3896
rect 207256 3884 207262 3936
rect 216858 3884 216864 3936
rect 216916 3924 216922 3936
rect 231946 3924 231952 3936
rect 216916 3896 231952 3924
rect 216916 3884 216922 3896
rect 231946 3884 231952 3896
rect 232004 3884 232010 3936
rect 252646 3884 252652 3936
rect 252704 3924 252710 3936
rect 265342 3924 265348 3936
rect 252704 3896 265348 3924
rect 252704 3884 252710 3896
rect 265342 3884 265348 3896
rect 265400 3884 265406 3936
rect 336734 3884 336740 3936
rect 336792 3924 336798 3936
rect 458082 3924 458088 3936
rect 336792 3896 458088 3924
rect 336792 3884 336798 3896
rect 458082 3884 458088 3896
rect 458140 3884 458146 3936
rect 160186 3816 160192 3868
rect 160244 3856 160250 3868
rect 205726 3856 205732 3868
rect 160244 3828 205732 3856
rect 160244 3816 160250 3828
rect 205726 3816 205732 3828
rect 205784 3816 205790 3868
rect 213362 3816 213368 3868
rect 213420 3856 213426 3868
rect 229186 3856 229192 3868
rect 213420 3828 229192 3856
rect 213420 3816 213426 3828
rect 229186 3816 229192 3828
rect 229244 3816 229250 3868
rect 252738 3816 252744 3868
rect 252796 3856 252802 3868
rect 266538 3856 266544 3868
rect 252796 3828 266544 3856
rect 252796 3816 252802 3828
rect 266538 3816 266544 3828
rect 266596 3816 266602 3868
rect 339494 3816 339500 3868
rect 339552 3856 339558 3868
rect 465166 3856 465172 3868
rect 339552 3828 465172 3856
rect 339552 3816 339558 3828
rect 465166 3816 465172 3828
rect 465224 3816 465230 3868
rect 574738 3816 574744 3868
rect 574796 3856 574802 3868
rect 577406 3856 577412 3868
rect 574796 3828 577412 3856
rect 574796 3816 574802 3828
rect 577406 3816 577412 3828
rect 577464 3816 577470 3868
rect 156690 3748 156696 3800
rect 156748 3788 156754 3800
rect 204254 3788 204260 3800
rect 156748 3760 204260 3788
rect 156748 3748 156754 3760
rect 204254 3748 204260 3760
rect 204312 3748 204318 3800
rect 212166 3748 212172 3800
rect 212224 3788 212230 3800
rect 229370 3788 229376 3800
rect 212224 3760 229376 3788
rect 212224 3748 212230 3760
rect 229370 3748 229376 3760
rect 229428 3748 229434 3800
rect 253934 3748 253940 3800
rect 253992 3788 253998 3800
rect 270034 3788 270040 3800
rect 253992 3760 270040 3788
rect 253992 3748 253998 3760
rect 270034 3748 270040 3760
rect 270092 3748 270098 3800
rect 340874 3748 340880 3800
rect 340932 3788 340938 3800
rect 468662 3788 468668 3800
rect 340932 3760 468668 3788
rect 340932 3748 340938 3760
rect 468662 3748 468668 3760
rect 468720 3748 468726 3800
rect 153010 3680 153016 3732
rect 153068 3720 153074 3732
rect 203058 3720 203064 3732
rect 153068 3692 203064 3720
rect 153068 3680 153074 3692
rect 203058 3680 203064 3692
rect 203116 3680 203122 3732
rect 209774 3680 209780 3732
rect 209832 3720 209838 3732
rect 209832 3692 223712 3720
rect 209832 3680 209838 3692
rect 149514 3612 149520 3664
rect 149572 3652 149578 3664
rect 201586 3652 201592 3664
rect 149572 3624 201592 3652
rect 149572 3612 149578 3624
rect 201586 3612 201592 3624
rect 201644 3612 201650 3664
rect 208578 3612 208584 3664
rect 208636 3652 208642 3664
rect 223684 3652 223712 3692
rect 227530 3680 227536 3732
rect 227588 3720 227594 3732
rect 236178 3720 236184 3732
rect 227588 3692 236184 3720
rect 227588 3680 227594 3692
rect 236178 3680 236184 3692
rect 236236 3680 236242 3732
rect 238110 3680 238116 3732
rect 238168 3720 238174 3732
rect 240318 3720 240324 3732
rect 238168 3692 240324 3720
rect 238168 3680 238174 3692
rect 240318 3680 240324 3692
rect 240376 3680 240382 3732
rect 255314 3680 255320 3732
rect 255372 3720 255378 3732
rect 273622 3720 273628 3732
rect 255372 3692 273628 3720
rect 255372 3680 255378 3692
rect 273622 3680 273628 3692
rect 273680 3680 273686 3732
rect 342254 3680 342260 3732
rect 342312 3720 342318 3732
rect 472250 3720 472256 3732
rect 342312 3692 472256 3720
rect 342312 3680 342318 3692
rect 472250 3680 472256 3692
rect 472308 3680 472314 3732
rect 227898 3652 227904 3664
rect 208636 3624 219434 3652
rect 223684 3624 227904 3652
rect 208636 3612 208642 3624
rect 145926 3544 145932 3596
rect 145984 3584 145990 3596
rect 200114 3584 200120 3596
rect 145984 3556 200120 3584
rect 145984 3544 145990 3556
rect 200114 3544 200120 3556
rect 200172 3544 200178 3596
rect 219406 3584 219434 3624
rect 227898 3612 227904 3624
rect 227956 3612 227962 3664
rect 229830 3612 229836 3664
rect 229888 3652 229894 3664
rect 237466 3652 237472 3664
rect 229888 3624 237472 3652
rect 229888 3612 229894 3624
rect 237466 3612 237472 3624
rect 237524 3612 237530 3664
rect 245654 3612 245660 3664
rect 245712 3652 245718 3664
rect 251174 3652 251180 3664
rect 245712 3624 251180 3652
rect 245712 3612 245718 3624
rect 251174 3612 251180 3624
rect 251232 3612 251238 3664
rect 258074 3612 258080 3664
rect 258132 3652 258138 3664
rect 277118 3652 277124 3664
rect 258132 3624 277124 3652
rect 258132 3612 258138 3624
rect 277118 3612 277124 3624
rect 277176 3612 277182 3664
rect 343634 3612 343640 3664
rect 343692 3652 343698 3664
rect 475746 3652 475752 3664
rect 343692 3624 475752 3652
rect 343692 3612 343698 3624
rect 475746 3612 475752 3624
rect 475804 3612 475810 3664
rect 227806 3584 227812 3596
rect 219406 3556 227812 3584
rect 227806 3544 227812 3556
rect 227864 3544 227870 3596
rect 232222 3544 232228 3596
rect 232280 3584 232286 3596
rect 235258 3584 235264 3596
rect 232280 3556 235264 3584
rect 232280 3544 232286 3556
rect 235258 3544 235264 3556
rect 235316 3544 235322 3596
rect 244366 3544 244372 3596
rect 244424 3584 244430 3596
rect 247586 3584 247592 3596
rect 244424 3556 247592 3584
rect 244424 3544 244430 3556
rect 247586 3544 247592 3556
rect 247644 3544 247650 3596
rect 249886 3544 249892 3596
rect 249944 3544 249950 3596
rect 251818 3544 251824 3596
rect 251876 3584 251882 3596
rect 254670 3584 254676 3596
rect 251876 3556 254676 3584
rect 251876 3544 251882 3556
rect 254670 3544 254676 3556
rect 254728 3544 254734 3596
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 280706 3584 280712 3596
rect 259512 3556 280712 3584
rect 259512 3544 259518 3556
rect 280706 3544 280712 3556
rect 280764 3544 280770 3596
rect 324406 3544 324412 3596
rect 324464 3584 324470 3596
rect 325602 3584 325608 3596
rect 324464 3556 325608 3584
rect 324464 3544 324470 3556
rect 325602 3544 325608 3556
rect 325660 3544 325666 3596
rect 332686 3544 332692 3596
rect 332744 3584 332750 3596
rect 333882 3584 333888 3596
rect 332744 3556 333888 3584
rect 332744 3544 332750 3556
rect 333882 3544 333888 3556
rect 333940 3544 333946 3596
rect 390646 3544 390652 3596
rect 390704 3584 390710 3596
rect 391842 3584 391848 3596
rect 390704 3556 391848 3584
rect 390704 3544 390710 3556
rect 391842 3544 391848 3556
rect 391900 3544 391906 3596
rect 391934 3544 391940 3596
rect 391992 3584 391998 3596
rect 582190 3584 582196 3596
rect 391992 3556 582196 3584
rect 391992 3544 391998 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 126974 3476 126980 3528
rect 127032 3516 127038 3528
rect 128998 3516 129004 3528
rect 127032 3488 129004 3516
rect 127032 3476 127038 3488
rect 128998 3476 129004 3488
rect 129056 3476 129062 3528
rect 134150 3476 134156 3528
rect 134208 3516 134214 3528
rect 137278 3516 137284 3528
rect 134208 3488 137284 3516
rect 134208 3476 134214 3488
rect 137278 3476 137284 3488
rect 137336 3476 137342 3528
rect 142430 3476 142436 3528
rect 142488 3516 142494 3528
rect 198734 3516 198740 3528
rect 142488 3488 198740 3516
rect 142488 3476 142494 3488
rect 198734 3476 198740 3488
rect 198792 3476 198798 3528
rect 199102 3476 199108 3528
rect 199160 3516 199166 3528
rect 223574 3516 223580 3528
rect 199160 3488 223580 3516
rect 199160 3476 199166 3488
rect 223574 3476 223580 3488
rect 223632 3476 223638 3528
rect 223942 3476 223948 3528
rect 224000 3516 224006 3528
rect 234614 3516 234620 3528
rect 224000 3488 234620 3516
rect 224000 3476 224006 3488
rect 234614 3476 234620 3488
rect 234672 3476 234678 3528
rect 239306 3476 239312 3528
rect 239364 3516 239370 3528
rect 240778 3516 240784 3528
rect 239364 3488 240784 3516
rect 239364 3476 239370 3488
rect 240778 3476 240784 3488
rect 240836 3476 240842 3528
rect 249904 3516 249932 3544
rect 258258 3516 258264 3528
rect 249904 3488 258264 3516
rect 258258 3476 258264 3488
rect 258316 3476 258322 3528
rect 260834 3476 260840 3528
rect 260892 3516 260898 3528
rect 284294 3516 284300 3528
rect 260892 3488 284300 3516
rect 260892 3476 260898 3488
rect 284294 3476 284300 3488
rect 284352 3476 284358 3528
rect 299566 3476 299572 3528
rect 299624 3516 299630 3528
rect 300762 3516 300768 3528
rect 299624 3488 300768 3516
rect 299624 3476 299630 3488
rect 300762 3476 300768 3488
rect 300820 3476 300826 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 316034 3476 316040 3528
rect 316092 3516 316098 3528
rect 317322 3516 317328 3528
rect 316092 3488 317328 3516
rect 316092 3476 316098 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 345014 3476 345020 3528
rect 345072 3516 345078 3528
rect 345072 3488 473216 3516
rect 345072 3476 345078 3488
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 193582 3448 193588 3460
rect 131816 3420 193588 3448
rect 131816 3408 131822 3420
rect 193582 3408 193588 3420
rect 193640 3408 193646 3460
rect 195606 3408 195612 3460
rect 195664 3448 195670 3460
rect 221090 3448 221096 3460
rect 195664 3420 221096 3448
rect 195664 3408 195670 3420
rect 221090 3408 221096 3420
rect 221148 3408 221154 3460
rect 231026 3408 231032 3460
rect 231084 3448 231090 3460
rect 237650 3448 237656 3460
rect 231084 3420 237656 3448
rect 231084 3408 231090 3420
rect 237650 3408 237656 3420
rect 237708 3408 237714 3460
rect 240502 3408 240508 3460
rect 240560 3448 240566 3460
rect 241790 3448 241796 3460
rect 240560 3420 241796 3448
rect 240560 3408 240566 3420
rect 241790 3408 241796 3420
rect 241848 3408 241854 3460
rect 250070 3408 250076 3460
rect 250128 3448 250134 3460
rect 259454 3448 259460 3460
rect 250128 3420 259460 3448
rect 250128 3408 250134 3420
rect 259454 3408 259460 3420
rect 259512 3408 259518 3460
rect 262398 3408 262404 3460
rect 262456 3448 262462 3460
rect 287790 3448 287796 3460
rect 262456 3420 287796 3448
rect 262456 3408 262462 3420
rect 287790 3408 287796 3420
rect 287848 3408 287854 3460
rect 365714 3408 365720 3460
rect 365772 3448 365778 3460
rect 367002 3448 367008 3460
rect 365772 3420 367008 3448
rect 365772 3408 365778 3420
rect 367002 3408 367008 3420
rect 367060 3408 367066 3460
rect 382274 3408 382280 3460
rect 382332 3448 382338 3460
rect 383562 3448 383568 3460
rect 382332 3420 383568 3448
rect 382332 3408 382338 3420
rect 383562 3408 383568 3420
rect 383620 3408 383626 3460
rect 391014 3408 391020 3460
rect 391072 3448 391078 3460
rect 391934 3448 391940 3460
rect 391072 3420 391940 3448
rect 391072 3408 391078 3420
rect 391934 3408 391940 3420
rect 391992 3408 391998 3460
rect 392026 3408 392032 3460
rect 392084 3448 392090 3460
rect 392084 3420 470594 3448
rect 392084 3408 392090 3420
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 141418 3380 141424 3392
rect 135312 3352 141424 3380
rect 135312 3340 135318 3352
rect 141418 3340 141424 3352
rect 141476 3340 141482 3392
rect 155402 3340 155408 3392
rect 155460 3380 155466 3392
rect 156598 3380 156604 3392
rect 155460 3352 156604 3380
rect 155460 3340 155466 3352
rect 156598 3340 156604 3352
rect 156656 3340 156662 3392
rect 160094 3340 160100 3392
rect 160152 3380 160158 3392
rect 161290 3380 161296 3392
rect 160152 3352 161296 3380
rect 160152 3340 160158 3352
rect 161290 3340 161296 3352
rect 161348 3340 161354 3392
rect 181438 3340 181444 3392
rect 181496 3380 181502 3392
rect 215294 3380 215300 3392
rect 181496 3352 215300 3380
rect 181496 3340 181502 3352
rect 215294 3340 215300 3352
rect 215352 3340 215358 3392
rect 222746 3340 222752 3392
rect 222804 3380 222810 3392
rect 233326 3380 233332 3392
rect 222804 3352 233332 3380
rect 222804 3340 222810 3352
rect 233326 3340 233332 3352
rect 233384 3340 233390 3392
rect 324314 3340 324320 3392
rect 324372 3380 324378 3392
rect 324372 3352 423720 3380
rect 324372 3340 324378 3352
rect 144730 3272 144736 3324
rect 144788 3312 144794 3324
rect 148318 3312 148324 3324
rect 144788 3284 148324 3312
rect 144788 3272 144794 3284
rect 148318 3272 148324 3284
rect 148376 3272 148382 3324
rect 188522 3272 188528 3324
rect 188580 3312 188586 3324
rect 218146 3312 218152 3324
rect 188580 3284 218152 3312
rect 188580 3272 188586 3284
rect 218146 3272 218152 3284
rect 218204 3272 218210 3324
rect 225138 3272 225144 3324
rect 225196 3312 225202 3324
rect 234798 3312 234804 3324
rect 225196 3284 234804 3312
rect 225196 3272 225202 3284
rect 234798 3272 234804 3284
rect 234856 3272 234862 3324
rect 248506 3272 248512 3324
rect 248564 3312 248570 3324
rect 257062 3312 257068 3324
rect 248564 3284 257068 3312
rect 248564 3272 248570 3284
rect 257062 3272 257068 3284
rect 257120 3272 257126 3324
rect 321554 3272 321560 3324
rect 321612 3312 321618 3324
rect 422570 3312 422576 3324
rect 321612 3284 422576 3312
rect 321612 3272 321618 3284
rect 422570 3272 422576 3284
rect 422628 3272 422634 3324
rect 423692 3312 423720 3352
rect 423766 3340 423772 3392
rect 423824 3380 423830 3392
rect 424962 3380 424968 3392
rect 423824 3352 424968 3380
rect 423824 3340 423830 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 431954 3340 431960 3392
rect 432012 3380 432018 3392
rect 433242 3380 433248 3392
rect 432012 3352 433248 3380
rect 432012 3340 432018 3352
rect 433242 3340 433248 3352
rect 433300 3340 433306 3392
rect 440326 3340 440332 3392
rect 440384 3380 440390 3392
rect 441522 3380 441528 3392
rect 440384 3352 441528 3380
rect 440384 3340 440390 3352
rect 441522 3340 441528 3352
rect 441580 3340 441586 3392
rect 429654 3312 429660 3324
rect 423692 3284 429660 3312
rect 429654 3272 429660 3284
rect 429712 3272 429718 3324
rect 470566 3312 470594 3420
rect 473188 3380 473216 3488
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474182 3516 474188 3528
rect 473412 3488 474188 3516
rect 473412 3476 473418 3488
rect 474182 3476 474188 3488
rect 474240 3476 474246 3528
rect 489914 3476 489920 3528
rect 489972 3516 489978 3528
rect 490742 3516 490748 3528
rect 489972 3488 490748 3516
rect 489972 3476 489978 3488
rect 490742 3476 490748 3488
rect 490800 3476 490806 3528
rect 498194 3476 498200 3528
rect 498252 3516 498258 3528
rect 499022 3516 499028 3528
rect 498252 3488 499028 3516
rect 498252 3476 498258 3488
rect 499022 3476 499028 3488
rect 499080 3476 499086 3528
rect 514754 3476 514760 3528
rect 514812 3516 514818 3528
rect 515582 3516 515588 3528
rect 514812 3488 515588 3516
rect 514812 3476 514818 3488
rect 515582 3476 515588 3488
rect 515640 3476 515646 3528
rect 523034 3476 523040 3528
rect 523092 3516 523098 3528
rect 523862 3516 523868 3528
rect 523092 3488 523868 3516
rect 523092 3476 523098 3488
rect 523862 3476 523868 3488
rect 523920 3476 523926 3528
rect 539594 3476 539600 3528
rect 539652 3516 539658 3528
rect 540422 3516 540428 3528
rect 539652 3488 540428 3516
rect 539652 3476 539658 3488
rect 540422 3476 540428 3488
rect 540480 3476 540486 3528
rect 564434 3476 564440 3528
rect 564492 3516 564498 3528
rect 565262 3516 565268 3528
rect 564492 3488 565268 3516
rect 564492 3476 564498 3488
rect 565262 3476 565268 3488
rect 565320 3476 565326 3528
rect 570598 3476 570604 3528
rect 570656 3516 570662 3528
rect 571518 3516 571524 3528
rect 570656 3488 571524 3516
rect 570656 3476 570662 3488
rect 571518 3476 571524 3488
rect 571576 3476 571582 3528
rect 580994 3448 581000 3460
rect 480226 3420 581000 3448
rect 479334 3380 479340 3392
rect 473188 3352 479340 3380
rect 479334 3340 479340 3352
rect 479392 3340 479398 3392
rect 480226 3312 480254 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 470566 3284 480254 3312
rect 192018 3204 192024 3256
rect 192076 3244 192082 3256
rect 219710 3244 219716 3256
rect 192076 3216 219716 3244
rect 192076 3204 192082 3216
rect 219710 3204 219716 3216
rect 219768 3204 219774 3256
rect 226334 3204 226340 3256
rect 226392 3244 226398 3256
rect 235994 3244 236000 3256
rect 226392 3216 236000 3244
rect 226392 3204 226398 3216
rect 235994 3204 236000 3216
rect 236052 3204 236058 3256
rect 317506 3204 317512 3256
rect 317564 3244 317570 3256
rect 415394 3244 415400 3256
rect 317564 3216 415400 3244
rect 317564 3204 317570 3216
rect 415394 3204 415400 3216
rect 415452 3204 415458 3256
rect 415486 3204 415492 3256
rect 415544 3244 415550 3256
rect 416682 3244 416688 3256
rect 415544 3216 416688 3244
rect 415544 3204 415550 3216
rect 416682 3204 416688 3216
rect 416740 3204 416746 3256
rect 151814 3136 151820 3188
rect 151872 3176 151878 3188
rect 155218 3176 155224 3188
rect 151872 3148 155224 3176
rect 151872 3136 151878 3148
rect 155218 3136 155224 3148
rect 155276 3136 155282 3188
rect 221550 3136 221556 3188
rect 221608 3176 221614 3188
rect 233602 3176 233608 3188
rect 221608 3148 233608 3176
rect 221608 3136 221614 3148
rect 233602 3136 233608 3148
rect 233660 3136 233666 3188
rect 390554 3136 390560 3188
rect 390612 3176 390618 3188
rect 392026 3176 392032 3188
rect 390612 3148 392032 3176
rect 390612 3136 390618 3148
rect 392026 3136 392032 3148
rect 392084 3136 392090 3188
rect 398926 3136 398932 3188
rect 398984 3176 398990 3188
rect 400122 3176 400128 3188
rect 398984 3148 400128 3176
rect 398984 3136 398990 3148
rect 400122 3136 400128 3148
rect 400180 3136 400186 3188
rect 407206 3136 407212 3188
rect 407264 3176 407270 3188
rect 408402 3176 408408 3188
rect 407264 3148 408408 3176
rect 407264 3136 407270 3148
rect 408402 3136 408408 3148
rect 408460 3136 408466 3188
rect 205082 3068 205088 3120
rect 205140 3108 205146 3120
rect 226518 3108 226524 3120
rect 205140 3080 226524 3108
rect 205140 3068 205146 3080
rect 226518 3068 226524 3080
rect 226576 3068 226582 3120
rect 137646 3000 137652 3052
rect 137704 3040 137710 3052
rect 140038 3040 140044 3052
rect 137704 3012 140044 3040
rect 137704 3000 137710 3012
rect 140038 3000 140044 3012
rect 140096 3000 140102 3052
rect 234614 3000 234620 3052
rect 234672 3040 234678 3052
rect 238938 3040 238944 3052
rect 234672 3012 238944 3040
rect 234672 3000 234678 3012
rect 238938 3000 238944 3012
rect 238996 3000 239002 3052
rect 248598 3000 248604 3052
rect 248656 3040 248662 3052
rect 255866 3040 255872 3052
rect 248656 3012 255872 3040
rect 248656 3000 248662 3012
rect 255866 3000 255872 3012
rect 255924 3000 255930 3052
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 573910 3040 573916 3052
rect 572036 3012 573916 3040
rect 572036 3000 572042 3012
rect 573910 3000 573916 3012
rect 573968 3000 573974 3052
rect 148318 2932 148324 2984
rect 148376 2972 148382 2984
rect 152458 2972 152464 2984
rect 148376 2944 152464 2972
rect 148376 2932 148382 2944
rect 152458 2932 152464 2944
rect 152516 2932 152522 2984
rect 233418 2864 233424 2916
rect 233476 2904 233482 2916
rect 238018 2904 238024 2916
rect 233476 2876 238024 2904
rect 233476 2864 233482 2876
rect 238018 2864 238024 2876
rect 238076 2864 238082 2916
rect 448514 1912 448520 1964
rect 448572 1952 448578 1964
rect 449802 1952 449808 1964
rect 448572 1924 449808 1952
rect 448572 1912 448578 1924
rect 449802 1912 449808 1924
rect 449860 1912 449866 1964
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 292580 700884 292632 700936
rect 332508 700884 332560 700936
rect 295340 700816 295392 700868
rect 348792 700816 348844 700868
rect 298100 700748 298152 700800
rect 364984 700748 365036 700800
rect 300860 700680 300912 700732
rect 397460 700680 397512 700732
rect 302240 700612 302292 700664
rect 413652 700612 413704 700664
rect 305000 700544 305052 700596
rect 429844 700544 429896 700596
rect 307760 700476 307812 700528
rect 462320 700476 462372 700528
rect 310520 700408 310572 700460
rect 478512 700408 478564 700460
rect 316040 700340 316092 700392
rect 527180 700340 527232 700392
rect 170312 700272 170364 700324
rect 192484 700272 192536 700324
rect 202788 700272 202840 700324
rect 220084 700272 220136 700324
rect 235172 700272 235224 700324
rect 282184 700272 282236 700324
rect 291844 700272 291896 700324
rect 300124 700272 300176 700324
rect 318800 700272 318852 700324
rect 543464 700272 543516 700324
rect 283840 700068 283892 700120
rect 284944 700068 284996 700120
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 322940 696940 322992 696992
rect 580172 696940 580224 696992
rect 3424 683136 3476 683188
rect 93124 683136 93176 683188
rect 325700 683136 325752 683188
rect 580172 683136 580224 683188
rect 328460 670692 328512 670744
rect 580172 670692 580224 670744
rect 3516 656888 3568 656940
rect 246304 656888 246356 656940
rect 331220 643084 331272 643136
rect 580172 643084 580224 643136
rect 3516 632068 3568 632120
rect 244280 632068 244332 632120
rect 333980 630640 334032 630692
rect 580172 630640 580224 630692
rect 336740 616836 336792 616888
rect 580172 616836 580224 616888
rect 3332 605820 3384 605872
rect 238024 605820 238076 605872
rect 338120 590656 338172 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 235264 579640 235316 579692
rect 340880 576852 340932 576904
rect 580172 576852 580224 576904
rect 343640 563048 343692 563100
rect 579804 563048 579856 563100
rect 346400 536800 346452 536852
rect 580172 536800 580224 536852
rect 2964 527144 3016 527196
rect 228364 527144 228416 527196
rect 349160 524424 349212 524476
rect 580172 524424 580224 524476
rect 3332 514768 3384 514820
rect 226340 514768 226392 514820
rect 351920 510620 351972 510672
rect 580172 510620 580224 510672
rect 354680 484372 354732 484424
rect 580172 484372 580224 484424
rect 220084 476756 220136 476808
rect 277400 476756 277452 476808
rect 2872 474716 2924 474768
rect 220084 474716 220136 474768
rect 356060 470568 356112 470620
rect 579988 470568 580040 470620
rect 358820 456764 358872 456816
rect 580172 456764 580224 456816
rect 361580 430584 361632 430636
rect 580172 430584 580224 430636
rect 2780 423512 2832 423564
rect 4804 423512 4856 423564
rect 364340 418140 364392 418192
rect 580172 418140 580224 418192
rect 3332 409844 3384 409896
rect 211160 409844 211212 409896
rect 367100 404336 367152 404388
rect 580172 404336 580224 404388
rect 369860 378156 369912 378208
rect 580172 378156 580224 378208
rect 136640 371832 136692 371884
rect 269672 371832 269724 371884
rect 3332 371220 3384 371272
rect 13820 371220 13872 371272
rect 93124 370472 93176 370524
rect 251824 370472 251876 370524
rect 13820 369112 13872 369164
rect 205640 369112 205692 369164
rect 4804 367752 4856 367804
rect 213184 367752 213236 367804
rect 40040 366324 40092 366376
rect 259828 366324 259880 366376
rect 104900 364964 104952 365016
rect 267556 364964 267608 365016
rect 372712 364352 372764 364404
rect 580172 364352 580224 364404
rect 192484 363604 192536 363656
rect 275192 363604 275244 363656
rect 228364 363196 228416 363248
rect 229100 363196 229152 363248
rect 238024 363196 238076 363248
rect 239312 363196 239364 363248
rect 220084 362924 220136 362976
rect 221372 362924 221424 362976
rect 235264 362924 235316 362976
rect 236736 362924 236788 362976
rect 246304 362924 246356 362976
rect 247040 362924 247092 362976
rect 71780 362856 71832 362908
rect 262404 362856 262456 362908
rect 284944 362856 284996 362908
rect 288072 362856 288124 362908
rect 4068 362788 4120 362840
rect 208584 362788 208636 362840
rect 218060 362788 218112 362840
rect 280344 362788 280396 362840
rect 3976 362720 4028 362772
rect 216220 362720 216272 362772
rect 3884 362652 3936 362704
rect 218796 362652 218848 362704
rect 3792 362584 3844 362636
rect 223948 362584 224000 362636
rect 3700 362516 3752 362568
rect 231676 362516 231728 362568
rect 3608 362448 3660 362500
rect 234160 362448 234212 362500
rect 23480 362380 23532 362432
rect 257252 362380 257304 362432
rect 3516 362312 3568 362364
rect 241888 362312 241940 362364
rect 3424 362244 3476 362296
rect 249616 362244 249668 362296
rect 313648 362244 313700 362296
rect 494060 362244 494112 362296
rect 6920 362176 6972 362228
rect 254676 362176 254728 362228
rect 266360 362176 266412 362228
rect 285496 362176 285548 362228
rect 321376 362176 321428 362228
rect 558920 362176 558972 362228
rect 88340 362108 88392 362160
rect 264980 362108 265032 362160
rect 153200 362040 153252 362092
rect 272708 362040 272760 362092
rect 382924 361904 382976 361956
rect 479524 361904 479576 361956
rect 282184 361836 282236 361888
rect 282920 361836 282972 361888
rect 290648 361836 290700 361888
rect 291844 361836 291896 361888
rect 388076 361836 388128 361888
rect 486424 361836 486476 361888
rect 385500 361768 385552 361820
rect 483664 361768 483716 361820
rect 377772 361700 377824 361752
rect 485044 361700 485096 361752
rect 375196 361632 375248 361684
rect 482284 361632 482336 361684
rect 380348 361564 380400 361616
rect 489184 361564 489236 361616
rect 186964 360476 187016 360528
rect 195704 360476 195756 360528
rect 4804 360408 4856 360460
rect 198280 360408 198332 360460
rect 191104 360340 191156 360392
rect 200856 360340 200908 360392
rect 191748 360272 191800 360324
rect 203432 360272 203484 360324
rect 188344 360204 188396 360256
rect 193220 360204 193272 360256
rect 390928 359388 390980 359440
rect 391848 359388 391900 359440
rect 391848 358776 391900 358828
rect 406384 358776 406436 358828
rect 3332 358708 3384 358760
rect 191748 358708 191800 358760
rect 482284 353200 482336 353252
rect 580172 353200 580224 353252
rect 3148 346332 3200 346384
rect 191104 346332 191156 346384
rect 3424 343612 3476 343664
rect 189080 343612 189132 343664
rect 7564 333956 7616 334008
rect 189080 333956 189132 334008
rect 485044 325592 485096 325644
rect 580172 325592 580224 325644
rect 22744 324300 22796 324352
rect 189080 324300 189132 324352
rect 2780 319812 2832 319864
rect 4804 319812 4856 319864
rect 394332 314712 394384 314764
rect 395344 314712 395396 314764
rect 489184 313216 489236 313268
rect 580172 313216 580224 313268
rect 3516 306280 3568 306332
rect 186964 306280 187016 306332
rect 4804 303628 4856 303680
rect 189080 303628 189132 303680
rect 394332 303628 394384 303680
rect 554044 303628 554096 303680
rect 479524 299412 479576 299464
rect 580172 299412 580224 299464
rect 3056 293904 3108 293956
rect 188344 293904 188396 293956
rect 394424 284520 394476 284572
rect 399484 284520 399536 284572
rect 14464 274660 14516 274712
rect 189080 274660 189132 274712
rect 394424 274660 394476 274712
rect 551284 274660 551336 274712
rect 483664 273164 483716 273216
rect 580172 273164 580224 273216
rect 3516 267656 3568 267708
rect 7564 267656 7616 267708
rect 486424 259360 486476 259412
rect 580172 259360 580224 259412
rect 3608 253920 3660 253972
rect 189080 253920 189132 253972
rect 406384 245556 406436 245608
rect 580172 245556 580224 245608
rect 393780 244536 393832 244588
rect 396724 244536 396776 244588
rect 7564 244264 7616 244316
rect 189080 244264 189132 244316
rect 3424 241408 3476 241460
rect 189724 241408 189776 241460
rect 394148 233180 394200 233232
rect 579988 233180 580040 233232
rect 3516 224952 3568 225004
rect 189080 224952 189132 225004
rect 394056 219376 394108 219428
rect 580172 219376 580224 219428
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 21364 213936 21416 213988
rect 189080 213936 189132 213988
rect 394056 213936 394108 213988
rect 457444 213936 457496 213988
rect 393964 206932 394016 206984
rect 579804 206932 579856 206984
rect 3056 202784 3108 202836
rect 190092 202784 190144 202836
rect 3424 194556 3476 194608
rect 189080 194556 189132 194608
rect 394608 193128 394660 193180
rect 580172 193128 580224 193180
rect 3148 188980 3200 189032
rect 22744 188980 22796 189032
rect 394608 184900 394660 184952
rect 576124 184900 576176 184952
rect 395344 179324 395396 179376
rect 580172 179324 580224 179376
rect 308220 177760 308272 177812
rect 338764 177760 338816 177812
rect 320088 177692 320140 177744
rect 418160 177692 418212 177744
rect 188344 177624 188396 177676
rect 203708 177624 203760 177676
rect 209320 177624 209372 177676
rect 224960 177624 225012 177676
rect 323216 177624 323268 177676
rect 425060 177624 425112 177676
rect 191104 177556 191156 177608
rect 211436 177556 211488 177608
rect 227904 177556 227956 177608
rect 236644 177556 236696 177608
rect 326528 177556 326580 177608
rect 431960 177556 432012 177608
rect 184940 177488 184992 177540
rect 217140 177488 217192 177540
rect 248236 177488 248288 177540
rect 251824 177488 251876 177540
rect 262220 177488 262272 177540
rect 265256 177488 265308 177540
rect 282184 177488 282236 177540
rect 290188 177488 290240 177540
rect 300032 177488 300084 177540
rect 300860 177488 300912 177540
rect 309968 177488 310020 177540
rect 329656 177488 329708 177540
rect 440240 177488 440292 177540
rect 176660 177420 176712 177472
rect 214012 177420 214064 177472
rect 214564 177420 214616 177472
rect 225788 177420 225840 177472
rect 248144 177420 248196 177472
rect 252560 177420 252612 177472
rect 285680 177420 285732 177472
rect 286232 177420 286284 177472
rect 307024 177420 307076 177472
rect 332508 177420 332560 177472
rect 447140 177420 447192 177472
rect 141424 177352 141476 177404
rect 195428 177352 195480 177404
rect 206284 177352 206336 177404
rect 226892 177352 226944 177404
rect 246212 177352 246264 177404
rect 250076 177352 250128 177404
rect 252192 177352 252244 177404
rect 262220 177352 262272 177404
rect 264520 177352 264572 177404
rect 291200 177352 291252 177404
rect 302148 177352 302200 177404
rect 312544 177352 312596 177404
rect 315948 177352 316000 177404
rect 320824 177352 320876 177404
rect 335360 177352 335412 177404
rect 454040 177352 454092 177404
rect 134524 177284 134576 177336
rect 192300 177284 192352 177336
rect 201500 177284 201552 177336
rect 225420 177284 225472 177336
rect 247592 177284 247644 177336
rect 251272 177284 251324 177336
rect 252376 177284 252428 177336
rect 263600 177284 263652 177336
rect 281724 177284 281776 177336
rect 329104 177284 329156 177336
rect 338488 177284 338540 177336
rect 460940 177284 460992 177336
rect 246120 177216 246172 177268
rect 248420 177216 248472 177268
rect 343640 177148 343692 177200
rect 346952 177148 347004 177200
rect 333152 177080 333204 177132
rect 336188 177080 336240 177132
rect 373724 177012 373776 177064
rect 374644 177012 374696 177064
rect 226340 176944 226392 176996
rect 229192 176944 229244 176996
rect 238024 176944 238076 176996
rect 238852 176944 238904 176996
rect 284208 176944 284260 176996
rect 287704 176944 287756 176996
rect 217600 176876 217652 176928
rect 221188 176876 221240 176928
rect 234712 176876 234764 176928
rect 240232 176876 240284 176928
rect 262128 176876 262180 176928
rect 269672 176876 269724 176928
rect 273168 176876 273220 176928
rect 278044 176876 278096 176928
rect 236276 176808 236328 176860
rect 240324 176808 240376 176860
rect 192484 176672 192536 176724
rect 193404 176672 193456 176724
rect 226984 176672 227036 176724
rect 227812 176672 227864 176724
rect 235264 176672 235316 176724
rect 238300 176672 238352 176724
rect 240784 176672 240836 176724
rect 241520 176672 241572 176724
rect 244832 176672 244884 176724
rect 245752 176672 245804 176724
rect 272984 176672 273036 176724
rect 273904 176672 273956 176724
rect 279056 176672 279108 176724
rect 282276 176672 282328 176724
rect 291016 176672 291068 176724
rect 295984 176672 296036 176724
rect 297456 176672 297508 176724
rect 304264 176672 304316 176724
rect 307576 176672 307628 176724
rect 309876 176672 309928 176724
rect 318892 176672 318944 176724
rect 323584 176672 323636 176724
rect 326988 176672 327040 176724
rect 329196 176672 329248 176724
rect 337476 176672 337528 176724
rect 338856 176672 338908 176724
rect 354956 176672 355008 176724
rect 359464 176672 359516 176724
rect 362868 176672 362920 176724
rect 363604 176672 363656 176724
rect 368848 176672 368900 176724
rect 371884 176672 371936 176724
rect 380716 176672 380768 176724
rect 381544 176672 381596 176724
rect 384488 176672 384540 176724
rect 385592 176672 385644 176724
rect 327356 176604 327408 176656
rect 327540 176604 327592 176656
rect 357716 176604 357768 176656
rect 357900 176604 357952 176656
rect 309600 175992 309652 176044
rect 394700 175992 394752 176044
rect 125600 175924 125652 175976
rect 223764 175924 223816 175976
rect 275928 175924 275980 175976
rect 316040 175924 316092 175976
rect 390376 175924 390428 175976
rect 579620 175924 579672 175976
rect 340972 175652 341024 175704
rect 341892 175652 341944 175704
rect 375380 175652 375432 175704
rect 376300 175652 376352 175704
rect 194600 175584 194652 175636
rect 194784 175584 194836 175636
rect 200212 175584 200264 175636
rect 201132 175584 201184 175636
rect 207204 175584 207256 175636
rect 207756 175584 207808 175636
rect 215300 175584 215352 175636
rect 215576 175584 215628 175636
rect 218060 175584 218112 175636
rect 218612 175584 218664 175636
rect 229192 175584 229244 175636
rect 230020 175584 230072 175636
rect 230480 175584 230532 175636
rect 230940 175584 230992 175636
rect 233332 175584 233384 175636
rect 234068 175584 234120 175636
rect 241704 175584 241756 175636
rect 242348 175584 242400 175636
rect 242900 175584 242952 175636
rect 243452 175584 243504 175636
rect 253940 175584 253992 175636
rect 254676 175584 254728 175636
rect 255320 175584 255372 175636
rect 256332 175584 256384 175636
rect 259552 175584 259604 175636
rect 260380 175584 260432 175636
rect 263692 175584 263744 175636
rect 264612 175584 264664 175636
rect 267832 175584 267884 175636
rect 268660 175584 268712 175636
rect 269120 175584 269172 175636
rect 269764 175584 269816 175636
rect 287060 175584 287112 175636
rect 287796 175584 287848 175636
rect 302332 175584 302384 175636
rect 303252 175584 303304 175636
rect 305184 175584 305236 175636
rect 305828 175584 305880 175636
rect 310520 175584 310572 175636
rect 311348 175584 311400 175636
rect 311900 175584 311952 175636
rect 312452 175584 312504 175636
rect 340880 175584 340932 175636
rect 341340 175584 341392 175636
rect 342260 175584 342312 175636
rect 342812 175584 342864 175636
rect 343640 175584 343692 175636
rect 344468 175584 344520 175636
rect 345020 175584 345072 175636
rect 345940 175584 345992 175636
rect 347780 175584 347832 175636
rect 348516 175584 348568 175636
rect 349160 175584 349212 175636
rect 350172 175584 350224 175636
rect 362960 175584 363012 175636
rect 363420 175584 363472 175636
rect 375472 175584 375524 175636
rect 375932 175584 375984 175636
rect 249800 175516 249852 175568
rect 250076 175516 250128 175568
rect 288440 175516 288492 175568
rect 289268 175516 289320 175568
rect 313372 175516 313424 175568
rect 313924 175516 313976 175568
rect 317512 175516 317564 175568
rect 318156 175516 318208 175568
rect 284300 175448 284352 175500
rect 284668 175448 284720 175500
rect 339500 175448 339552 175500
rect 339868 175448 339920 175500
rect 374000 175448 374052 175500
rect 374828 175448 374880 175500
rect 160100 174564 160152 174616
rect 207020 174564 207072 174616
rect 348424 174564 348476 174616
rect 483020 174564 483072 174616
rect 155224 174496 155276 174548
rect 202880 174496 202932 174548
rect 283656 174496 283708 174548
rect 333980 174496 334032 174548
rect 387708 174496 387760 174548
rect 571984 174496 572036 174548
rect 258264 174088 258316 174140
rect 258908 174088 258960 174140
rect 236092 173952 236144 174004
rect 236276 173952 236328 174004
rect 346400 173816 346452 173868
rect 347044 173816 347096 173868
rect 164240 173204 164292 173256
rect 208400 173204 208452 173256
rect 333336 173204 333388 173256
rect 448520 173204 448572 173256
rect 158720 173136 158772 173188
rect 205640 173136 205692 173188
rect 279148 173136 279200 173188
rect 324412 173136 324464 173188
rect 351736 173136 351788 173188
rect 489920 173136 489972 173188
rect 209964 171980 210016 172032
rect 226340 171980 226392 172032
rect 168380 171844 168432 171896
rect 209780 171844 209832 171896
rect 314752 171844 314804 171896
rect 407120 171844 407172 171896
rect 142804 171776 142856 171828
rect 198004 171776 198056 171828
rect 248512 171776 248564 171828
rect 248972 171776 249024 171828
rect 273260 171776 273312 171828
rect 273812 171776 273864 171828
rect 280160 171776 280212 171828
rect 280436 171776 280488 171828
rect 292580 171776 292632 171828
rect 293316 171776 293368 171828
rect 298100 171776 298152 171828
rect 299020 171776 299072 171828
rect 299480 171776 299532 171828
rect 300124 171776 300176 171828
rect 322940 171776 322992 171828
rect 323860 171776 323912 171828
rect 327172 171776 327224 171828
rect 327908 171776 327960 171828
rect 353300 171776 353352 171828
rect 353668 171776 353720 171828
rect 356152 171776 356204 171828
rect 356796 171776 356848 171828
rect 357440 171776 357492 171828
rect 358268 171776 358320 171828
rect 353392 171708 353444 171760
rect 354220 171708 354272 171760
rect 353208 171640 353260 171692
rect 494060 171776 494112 171828
rect 379520 171708 379572 171760
rect 379980 171708 380032 171760
rect 380900 171708 380952 171760
rect 381452 171708 381504 171760
rect 385040 171708 385092 171760
rect 385684 171708 385736 171760
rect 387800 171708 387852 171760
rect 388260 171708 388312 171760
rect 383660 171640 383712 171692
rect 384580 171640 384632 171692
rect 204260 171232 204312 171284
rect 204812 171232 204864 171284
rect 321652 171096 321704 171148
rect 322204 171096 322256 171148
rect 329932 171096 329984 171148
rect 330484 171096 330536 171148
rect 186320 170416 186372 170468
rect 218152 170416 218204 170468
rect 143540 170348 143592 170400
rect 198924 170348 198976 170400
rect 292764 170348 292816 170400
rect 356060 170348 356112 170400
rect 356336 170348 356388 170400
rect 500960 170348 501012 170400
rect 190460 169056 190512 169108
rect 219624 169056 219676 169108
rect 337660 169056 337712 169108
rect 459560 169056 459612 169108
rect 146300 168988 146352 169040
rect 200580 168988 200632 169040
rect 298192 168988 298244 169040
rect 298376 168988 298428 169040
rect 358912 168988 358964 169040
rect 507860 168988 507912 169040
rect 150440 167628 150492 167680
rect 202144 167628 202196 167680
rect 361856 167628 361908 167680
rect 514760 167628 514812 167680
rect 276112 167016 276164 167068
rect 276940 167016 276992 167068
rect 554044 166948 554096 167000
rect 580172 166948 580224 167000
rect 297548 166336 297600 166388
rect 367192 166336 367244 166388
rect 157340 166268 157392 166320
rect 205180 166268 205232 166320
rect 366456 166268 366508 166320
rect 525800 166268 525852 166320
rect 311992 164908 312044 164960
rect 400220 164908 400272 164960
rect 161480 164840 161532 164892
rect 207296 164840 207348 164892
rect 368480 164840 368532 164892
rect 529940 164840 529992 164892
rect 3332 164160 3384 164212
rect 14464 164160 14516 164212
rect 308312 163548 308364 163600
rect 391940 163548 391992 163600
rect 165620 163480 165672 163532
rect 208492 163480 208544 163532
rect 372804 163480 372856 163532
rect 539600 163480 539652 163532
rect 319076 162188 319128 162240
rect 416780 162188 416832 162240
rect 172520 162120 172572 162172
rect 211896 162120 211948 162172
rect 374184 162120 374236 162172
rect 543740 162120 543792 162172
rect 316224 160760 316276 160812
rect 411260 160760 411312 160812
rect 176752 160692 176804 160744
rect 212724 160692 212776 160744
rect 375472 160692 375524 160744
rect 547880 160692 547932 160744
rect 328460 159400 328512 159452
rect 438860 159400 438912 159452
rect 179420 159332 179472 159384
rect 215484 159332 215536 159384
rect 378416 159332 378468 159384
rect 554780 159332 554832 159384
rect 327264 158040 327316 158092
rect 434720 158040 434772 158092
rect 183560 157972 183612 158024
rect 216772 157972 216824 158024
rect 381544 157972 381596 158024
rect 557540 157972 557592 158024
rect 314660 156680 314712 156732
rect 407212 156680 407264 156732
rect 129740 156612 129792 156664
rect 192484 156612 192536 156664
rect 382188 156612 382240 156664
rect 561680 156612 561732 156664
rect 313464 155252 313516 155304
rect 404360 155252 404412 155304
rect 137284 155184 137336 155236
rect 194692 155184 194744 155236
rect 383752 155184 383804 155236
rect 564440 155184 564492 155236
rect 309232 153892 309284 153944
rect 396080 153892 396132 153944
rect 140044 153824 140096 153876
rect 196072 153824 196124 153876
rect 385132 153824 385184 153876
rect 568580 153824 568632 153876
rect 394516 153144 394568 153196
rect 580172 153144 580224 153196
rect 148324 152464 148376 152516
rect 199016 152464 199068 152516
rect 306472 152464 306524 152516
rect 389180 152464 389232 152516
rect 152464 151036 152516 151088
rect 200212 151036 200264 151088
rect 386604 151036 386656 151088
rect 572812 151036 572864 151088
rect 3332 150356 3384 150408
rect 190184 150356 190236 150408
rect 310796 149744 310848 149796
rect 398840 149744 398892 149796
rect 379612 149676 379664 149728
rect 556160 149676 556212 149728
rect 321744 148384 321796 148436
rect 423680 148384 423732 148436
rect 156604 148316 156656 148368
rect 204352 148316 204404 148368
rect 387984 148316 388036 148368
rect 574744 148316 574796 148368
rect 324504 146956 324556 147008
rect 430580 146956 430632 147008
rect 367284 146888 367336 146940
rect 528560 146888 528612 146940
rect 329840 145528 329892 145580
rect 440332 145528 440384 145580
rect 336004 144168 336056 144220
rect 448612 144168 448664 144220
rect 338856 142808 338908 142860
rect 458180 142808 458232 142860
rect 347780 141380 347832 141432
rect 484400 141380 484452 141432
rect 353484 140020 353536 140072
rect 495440 140020 495492 140072
rect 399484 139340 399536 139392
rect 579896 139340 579948 139392
rect 3056 137912 3108 137964
rect 190000 137912 190052 137964
rect 356244 137232 356296 137284
rect 502340 137232 502392 137284
rect 357532 135872 357584 135924
rect 506480 135872 506532 135924
rect 360384 134512 360436 134564
rect 513380 134512 513432 134564
rect 363604 133152 363656 133204
rect 516140 133152 516192 133204
rect 364340 131724 364392 131776
rect 520280 131724 520332 131776
rect 374644 130364 374696 130416
rect 540980 130364 541032 130416
rect 305276 129004 305328 129056
rect 385132 129004 385184 129056
rect 385684 129004 385736 129056
rect 565820 129004 565872 129056
rect 312544 127576 312596 127628
rect 376852 127576 376904 127628
rect 380992 127576 381044 127628
rect 558920 127576 558972 127628
rect 551284 126896 551336 126948
rect 579988 126896 580040 126948
rect 376944 126216 376996 126268
rect 550640 126216 550692 126268
rect 325700 124856 325752 124908
rect 432052 124856 432104 124908
rect 280436 123428 280488 123480
rect 329840 123428 329892 123480
rect 330024 123428 330076 123480
rect 441620 123428 441672 123480
rect 331404 122068 331456 122120
rect 445760 122068 445812 122120
rect 334164 120708 334216 120760
rect 452660 120708 452712 120760
rect 339592 119348 339644 119400
rect 463700 119348 463752 119400
rect 343824 117920 343876 117972
rect 473360 117920 473412 117972
rect 347872 116628 347924 116680
rect 288624 116560 288676 116612
rect 347780 116560 347832 116612
rect 481640 116560 481692 116612
rect 350540 115200 350592 115252
rect 490012 115200 490064 115252
rect 354680 113772 354732 113824
rect 499580 113772 499632 113824
rect 394424 113092 394476 113144
rect 580172 113092 580224 113144
rect 361580 111052 361632 111104
rect 514852 111052 514904 111104
rect 3332 110848 3384 110900
rect 7564 110848 7616 110900
rect 365812 109692 365864 109744
rect 524420 109692 524472 109744
rect 370136 108264 370188 108316
rect 535460 108264 535512 108316
rect 372620 106904 372672 106956
rect 539692 106904 539744 106956
rect 374092 105544 374144 105596
rect 542360 105544 542412 105596
rect 300860 104116 300912 104168
rect 375472 104116 375524 104168
rect 375564 104116 375616 104168
rect 546500 104116 546552 104168
rect 378324 102756 378376 102808
rect 553400 102756 553452 102808
rect 379520 101396 379572 101448
rect 556252 101396 556304 101448
rect 394332 100648 394384 100700
rect 580172 100648 580224 100700
rect 386420 98608 386472 98660
rect 570604 98608 570656 98660
rect 389272 97248 389324 97300
rect 578240 97248 578292 97300
rect 334072 94460 334124 94512
rect 451280 94460 451332 94512
rect 327172 93100 327224 93152
rect 437480 93100 437532 93152
rect 292764 91740 292816 91792
rect 357532 91740 357584 91792
rect 357624 91740 357676 91792
rect 505100 91740 505152 91792
rect 396724 86912 396776 86964
rect 580172 86912 580224 86964
rect 3332 85484 3384 85536
rect 189908 85484 189960 85536
rect 394240 73108 394292 73160
rect 580172 73108 580224 73160
rect 3332 71680 3384 71732
rect 21364 71680 21416 71732
rect 309140 61344 309192 61396
rect 393320 61344 393372 61396
rect 394148 60664 394200 60716
rect 580172 60664 580224 60716
rect 303712 59984 303764 60036
rect 382372 59984 382424 60036
rect 305184 58624 305236 58676
rect 386420 58624 386472 58676
rect 302424 57196 302476 57248
rect 379520 57196 379572 57248
rect 299572 55836 299624 55888
rect 372620 55836 372672 55888
rect 291384 54476 291436 54528
rect 354680 54476 354732 54528
rect 296720 53048 296772 53100
rect 365812 53048 365864 53100
rect 294144 51688 294196 51740
rect 361580 51688 361632 51740
rect 383660 51688 383712 51740
rect 566464 51688 566516 51740
rect 289820 50328 289872 50380
rect 350540 50328 350592 50380
rect 295984 48968 296036 49020
rect 352104 48968 352156 49020
rect 387892 48968 387944 49020
rect 574100 48968 574152 49020
rect 292580 47676 292632 47728
rect 357624 47676 357676 47728
rect 357440 47540 357492 47592
rect 506572 47540 506624 47592
rect 457444 46860 457496 46912
rect 580172 46860 580224 46912
rect 278872 46180 278924 46232
rect 325700 46180 325752 46232
rect 335544 46180 335596 46232
rect 456892 46180 456944 46232
rect 3516 45500 3568 45552
rect 189816 45500 189868 45552
rect 309876 44820 309928 44872
rect 374092 44820 374144 44872
rect 380900 44820 380952 44872
rect 560300 44820 560352 44872
rect 320824 43392 320876 43444
rect 408500 43392 408552 43444
rect 303620 42168 303672 42220
rect 382556 42168 382608 42220
rect 382464 42032 382516 42084
rect 564532 42032 564584 42084
rect 277492 40672 277544 40724
rect 323124 40672 323176 40724
rect 371884 40672 371936 40724
rect 531320 40672 531372 40724
rect 276296 39312 276348 39364
rect 318800 39312 318852 39364
rect 365720 39312 365772 39364
rect 523040 39312 523092 39364
rect 273352 37884 273404 37936
rect 311992 37884 312044 37936
rect 358820 37884 358872 37936
rect 509240 37884 509292 37936
rect 300124 36524 300176 36576
rect 349344 36524 349396 36576
rect 351920 36524 351972 36576
rect 491300 36524 491352 36576
rect 271880 35164 271932 35216
rect 307760 35164 307812 35216
rect 323032 35164 323084 35216
rect 426440 35164 426492 35216
rect 287704 33736 287756 33788
rect 335452 33736 335504 33788
rect 347044 33736 347096 33788
rect 473452 33736 473504 33788
rect 2872 33056 2924 33108
rect 190092 33056 190144 33108
rect 394056 33056 394108 33108
rect 579896 33056 579948 33108
rect 278044 32444 278096 32496
rect 310704 32444 310756 32496
rect 298284 32376 298336 32428
rect 368480 32376 368532 32428
rect 270500 31016 270552 31068
rect 305092 31016 305144 31068
rect 329196 31016 329248 31068
rect 433340 31016 433392 31068
rect 254124 29588 254176 29640
rect 267924 29588 267976 29640
rect 268016 29588 268068 29640
rect 299572 29588 299624 29640
rect 323584 29588 323636 29640
rect 415492 29588 415544 29640
rect 282276 28228 282328 28280
rect 324504 28228 324556 28280
rect 331220 28228 331272 28280
rect 444380 28228 444432 28280
rect 306380 26936 306432 26988
rect 387892 26936 387944 26988
rect 267832 26868 267884 26920
rect 300860 26868 300912 26920
rect 376760 26868 376812 26920
rect 549260 26868 549312 26920
rect 266544 25508 266596 25560
rect 298284 25508 298336 25560
rect 305000 25508 305052 25560
rect 383660 25508 383712 25560
rect 385040 25508 385092 25560
rect 569960 25508 570012 25560
rect 264980 24080 265032 24132
rect 294144 24080 294196 24132
rect 302332 24080 302384 24132
rect 380900 24080 380952 24132
rect 382280 24080 382332 24132
rect 563060 24080 563112 24132
rect 298192 22788 298244 22840
rect 370044 22788 370096 22840
rect 267740 22720 267792 22772
rect 299664 22720 299716 22772
rect 359464 22720 359516 22772
rect 498200 22720 498252 22772
rect 270684 21428 270736 21480
rect 307852 21428 307904 21480
rect 284392 21360 284444 21412
rect 336832 21360 336884 21412
rect 353392 21360 353444 21412
rect 498292 21360 498344 21412
rect 393964 20612 394016 20664
rect 579896 20612 579948 20664
rect 280252 20000 280304 20052
rect 327172 20000 327224 20052
rect 310612 19932 310664 19984
rect 397460 19932 397512 19984
rect 256792 18776 256844 18828
rect 276204 18776 276256 18828
rect 276112 18640 276164 18692
rect 320364 18640 320416 18692
rect 338764 18640 338816 18692
rect 390652 18640 390704 18692
rect 287152 18572 287204 18624
rect 343732 18572 343784 18624
rect 368572 18572 368624 18624
rect 531412 18572 531464 18624
rect 304264 17280 304316 17332
rect 365720 17280 365772 17332
rect 266360 17212 266412 17264
rect 295524 17212 295576 17264
rect 364524 17212 364576 17264
rect 523132 17212 523184 17264
rect 273904 15920 273956 15972
rect 309692 15920 309744 15972
rect 282920 15852 282972 15904
rect 332692 15852 332744 15904
rect 349436 15852 349488 15904
rect 487160 15852 487212 15904
rect 270592 14492 270644 14544
rect 306380 14492 306432 14544
rect 309784 14492 309836 14544
rect 390928 14492 390980 14544
rect 274732 14424 274784 14476
rect 316224 14424 316276 14476
rect 346492 14424 346544 14476
rect 480536 14424 480588 14476
rect 356152 13268 356204 13320
rect 503720 13268 503772 13320
rect 340972 13200 341024 13252
rect 341156 13200 341208 13252
rect 360200 13200 360252 13252
rect 511264 13200 511316 13252
rect 266452 13132 266504 13184
rect 297272 13132 297324 13184
rect 363052 13132 363104 13184
rect 517888 13132 517940 13184
rect 197912 13064 197964 13116
rect 222292 13064 222344 13116
rect 254032 13064 254084 13116
rect 267740 13064 267792 13116
rect 269212 13064 269264 13116
rect 303160 13064 303212 13116
rect 307024 13064 307076 13116
rect 340972 13064 341024 13116
rect 364432 13064 364484 13116
rect 521660 13064 521712 13116
rect 341064 12044 341116 12096
rect 467472 12044 467524 12096
rect 342352 11976 342404 12028
rect 470600 11976 470652 12028
rect 345204 11908 345256 11960
rect 478144 11908 478196 11960
rect 259644 11840 259696 11892
rect 281632 11840 281684 11892
rect 349252 11840 349304 11892
rect 486424 11840 486476 11892
rect 176660 11772 176712 11824
rect 177856 11772 177908 11824
rect 201500 11772 201552 11824
rect 202696 11772 202748 11824
rect 273260 11772 273312 11824
rect 313832 11772 313884 11824
rect 352012 11772 352064 11824
rect 493048 11772 493100 11824
rect 169576 11704 169628 11756
rect 209872 11704 209924 11756
rect 242900 11704 242952 11756
rect 244096 11704 244148 11756
rect 281540 11704 281592 11756
rect 329104 11704 329156 11756
rect 331220 11704 331272 11756
rect 353300 11704 353352 11756
rect 497096 11704 497148 11756
rect 332784 11636 332836 11688
rect 310520 10684 310572 10736
rect 398932 10684 398984 10736
rect 313280 10616 313332 10668
rect 403624 10616 403676 10668
rect 316132 10548 316184 10600
rect 410800 10548 410852 10600
rect 201684 10480 201736 10532
rect 209044 10480 209096 10532
rect 317604 10480 317656 10532
rect 414296 10480 414348 10532
rect 262496 10412 262548 10464
rect 288992 10412 289044 10464
rect 320272 10412 320324 10464
rect 420920 10412 420972 10464
rect 263784 10344 263836 10396
rect 289820 10344 289872 10396
rect 321652 10344 321704 10396
rect 423772 10344 423824 10396
rect 129004 10276 129056 10328
rect 191932 10276 191984 10328
rect 207112 10276 207164 10328
rect 226984 10276 227036 10328
rect 274640 10276 274692 10328
rect 314660 10276 314712 10328
rect 322940 10276 322992 10328
rect 428464 10276 428516 10328
rect 302240 9324 302292 9376
rect 378876 9324 378928 9376
rect 367100 9256 367152 9308
rect 527824 9256 527876 9308
rect 369952 9188 370004 9240
rect 534908 9188 534960 9240
rect 291292 9120 291344 9172
rect 354036 9120 354088 9172
rect 371332 9120 371384 9172
rect 538404 9120 538456 9172
rect 294052 9052 294104 9104
rect 361120 9052 361172 9104
rect 374000 9052 374052 9104
rect 545488 9052 545540 9104
rect 258356 8984 258408 9036
rect 278320 8984 278372 9036
rect 282184 8984 282236 9036
rect 293684 8984 293736 9036
rect 295432 8984 295484 9036
rect 364616 8984 364668 9036
rect 375380 8984 375432 9036
rect 549076 8984 549128 9036
rect 154212 8916 154264 8968
rect 188344 8916 188396 8968
rect 200304 8916 200356 8968
rect 223672 8916 223724 8968
rect 263692 8916 263744 8968
rect 292580 8916 292632 8968
rect 298100 8916 298152 8968
rect 371700 8916 371752 8968
rect 378140 8916 378192 8968
rect 552664 8916 552716 8968
rect 288532 8032 288584 8084
rect 346952 8032 347004 8084
rect 335360 7964 335412 8016
rect 455696 7964 455748 8016
rect 338120 7896 338172 7948
rect 462780 7896 462832 7948
rect 339684 7828 339736 7880
rect 466276 7828 466328 7880
rect 341156 7760 341208 7812
rect 469864 7760 469916 7812
rect 345112 7692 345164 7744
rect 476948 7692 477000 7744
rect 194416 7624 194468 7676
rect 217324 7624 217376 7676
rect 256700 7624 256752 7676
rect 274824 7624 274876 7676
rect 284484 7624 284536 7676
rect 339868 7624 339920 7676
rect 346400 7624 346452 7676
rect 481732 7624 481784 7676
rect 171968 7556 172020 7608
rect 191104 7556 191156 7608
rect 196808 7556 196860 7608
rect 222200 7556 222252 7608
rect 259552 7556 259604 7608
rect 283104 7556 283156 7608
rect 285864 7556 285916 7608
rect 343364 7556 343416 7608
rect 349160 7556 349212 7608
rect 488816 7556 488868 7608
rect 374092 7488 374144 7540
rect 375288 7488 375340 7540
rect 3424 6808 3476 6860
rect 189724 6808 189776 6860
rect 576124 6808 576176 6860
rect 580172 6808 580224 6860
rect 276112 6536 276164 6588
rect 318524 6536 318576 6588
rect 277400 6468 277452 6520
rect 322112 6468 322164 6520
rect 311900 6400 311952 6452
rect 402520 6400 402572 6452
rect 313372 6332 313424 6384
rect 406016 6332 406068 6384
rect 203892 6264 203944 6316
rect 214564 6264 214616 6316
rect 317420 6264 317472 6316
rect 413100 6264 413152 6316
rect 214472 6196 214524 6248
rect 230572 6196 230624 6248
rect 250076 6196 250128 6248
rect 260656 6196 260708 6248
rect 269120 6196 269172 6248
rect 304356 6196 304408 6248
rect 320180 6196 320232 6248
rect 420184 6196 420236 6248
rect 186136 6128 186188 6180
rect 216956 6128 217008 6180
rect 255504 6128 255556 6180
rect 272432 6128 272484 6180
rect 280160 6128 280212 6180
rect 329196 6128 329248 6180
rect 387800 6128 387852 6180
rect 576308 6128 576360 6180
rect 189724 5244 189776 5296
rect 219532 5244 219584 5296
rect 182548 5176 182600 5228
rect 215576 5176 215628 5228
rect 284300 5176 284352 5228
rect 338672 5176 338724 5228
rect 390744 5176 390796 5228
rect 391020 5176 391072 5228
rect 179052 5108 179104 5160
rect 214104 5108 214156 5160
rect 285772 5108 285824 5160
rect 342168 5108 342220 5160
rect 175464 5040 175516 5092
rect 212632 5040 212684 5092
rect 299480 5040 299532 5092
rect 374000 5040 374052 5092
rect 140136 4972 140188 5024
rect 197452 4972 197504 5024
rect 287060 4972 287112 5024
rect 345756 4972 345808 5024
rect 360292 4972 360344 5024
rect 512460 4972 512512 5024
rect 136456 4904 136508 4956
rect 195980 4904 196032 4956
rect 269764 4904 269816 4956
rect 285404 4904 285456 4956
rect 288440 4904 288492 4956
rect 349252 4904 349304 4956
rect 362960 4904 363012 4956
rect 519544 4972 519596 5024
rect 132960 4836 133012 4888
rect 194784 4836 194836 4888
rect 218060 4836 218112 4888
rect 232044 4836 232096 4888
rect 255412 4836 255464 4888
rect 271236 4836 271288 4888
rect 293960 4836 294012 4888
rect 359924 4836 359976 4888
rect 369860 4836 369912 4888
rect 533712 4836 533764 4888
rect 129372 4768 129424 4820
rect 193312 4768 193364 4820
rect 193220 4700 193272 4752
rect 220912 4768 220964 4820
rect 258264 4768 258316 4820
rect 279516 4768 279568 4820
rect 295340 4768 295392 4820
rect 363512 4768 363564 4820
rect 371240 4768 371292 4820
rect 537208 4768 537260 4820
rect 141240 4088 141292 4140
rect 142804 4088 142856 4140
rect 174268 4088 174320 4140
rect 212540 4088 212592 4140
rect 219256 4088 219308 4140
rect 232136 4088 232188 4140
rect 251180 4088 251232 4140
rect 261760 4088 261812 4140
rect 327080 4088 327132 4140
rect 436744 4088 436796 4140
rect 566464 4088 566516 4140
rect 568028 4088 568080 4140
rect 128176 4020 128228 4072
rect 134524 4020 134576 4072
rect 167184 4020 167236 4072
rect 208584 4020 208636 4072
rect 220452 4020 220504 4072
rect 233240 4020 233292 4072
rect 329932 4020 329984 4072
rect 443828 4020 443880 4072
rect 170772 3952 170824 4004
rect 211344 3952 211396 4004
rect 215668 3952 215720 4004
rect 230480 3952 230532 4004
rect 332600 3952 332652 4004
rect 450912 3952 450964 4004
rect 163688 3884 163740 3936
rect 207204 3884 207256 3936
rect 216864 3884 216916 3936
rect 231952 3884 232004 3936
rect 252652 3884 252704 3936
rect 265348 3884 265400 3936
rect 336740 3884 336792 3936
rect 458088 3884 458140 3936
rect 160192 3816 160244 3868
rect 205732 3816 205784 3868
rect 213368 3816 213420 3868
rect 229192 3816 229244 3868
rect 252744 3816 252796 3868
rect 266544 3816 266596 3868
rect 339500 3816 339552 3868
rect 465172 3816 465224 3868
rect 574744 3816 574796 3868
rect 577412 3816 577464 3868
rect 156696 3748 156748 3800
rect 204260 3748 204312 3800
rect 212172 3748 212224 3800
rect 229376 3748 229428 3800
rect 253940 3748 253992 3800
rect 270040 3748 270092 3800
rect 340880 3748 340932 3800
rect 468668 3748 468720 3800
rect 153016 3680 153068 3732
rect 203064 3680 203116 3732
rect 209780 3680 209832 3732
rect 149520 3612 149572 3664
rect 201592 3612 201644 3664
rect 208584 3612 208636 3664
rect 227536 3680 227588 3732
rect 236184 3680 236236 3732
rect 238116 3680 238168 3732
rect 240324 3680 240376 3732
rect 255320 3680 255372 3732
rect 273628 3680 273680 3732
rect 342260 3680 342312 3732
rect 472256 3680 472308 3732
rect 145932 3544 145984 3596
rect 200120 3544 200172 3596
rect 227904 3612 227956 3664
rect 229836 3612 229888 3664
rect 237472 3612 237524 3664
rect 245660 3612 245712 3664
rect 251180 3612 251232 3664
rect 258080 3612 258132 3664
rect 277124 3612 277176 3664
rect 343640 3612 343692 3664
rect 475752 3612 475804 3664
rect 227812 3544 227864 3596
rect 232228 3544 232280 3596
rect 235264 3544 235316 3596
rect 244372 3544 244424 3596
rect 247592 3544 247644 3596
rect 249892 3544 249944 3596
rect 251824 3544 251876 3596
rect 254676 3544 254728 3596
rect 259460 3544 259512 3596
rect 280712 3544 280764 3596
rect 324412 3544 324464 3596
rect 325608 3544 325660 3596
rect 332692 3544 332744 3596
rect 333888 3544 333940 3596
rect 390652 3544 390704 3596
rect 391848 3544 391900 3596
rect 391940 3544 391992 3596
rect 582196 3544 582248 3596
rect 126980 3476 127032 3528
rect 129004 3476 129056 3528
rect 134156 3476 134208 3528
rect 137284 3476 137336 3528
rect 142436 3476 142488 3528
rect 198740 3476 198792 3528
rect 199108 3476 199160 3528
rect 223580 3476 223632 3528
rect 223948 3476 224000 3528
rect 234620 3476 234672 3528
rect 239312 3476 239364 3528
rect 240784 3476 240836 3528
rect 258264 3476 258316 3528
rect 260840 3476 260892 3528
rect 284300 3476 284352 3528
rect 299572 3476 299624 3528
rect 300768 3476 300820 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 316040 3476 316092 3528
rect 317328 3476 317380 3528
rect 345020 3476 345072 3528
rect 131764 3408 131816 3460
rect 193588 3408 193640 3460
rect 195612 3408 195664 3460
rect 221096 3408 221148 3460
rect 231032 3408 231084 3460
rect 237656 3408 237708 3460
rect 240508 3408 240560 3460
rect 241796 3408 241848 3460
rect 250076 3408 250128 3460
rect 259460 3408 259512 3460
rect 262404 3408 262456 3460
rect 287796 3408 287848 3460
rect 365720 3408 365772 3460
rect 367008 3408 367060 3460
rect 382280 3408 382332 3460
rect 383568 3408 383620 3460
rect 391020 3408 391072 3460
rect 391940 3408 391992 3460
rect 392032 3408 392084 3460
rect 135260 3340 135312 3392
rect 141424 3340 141476 3392
rect 155408 3340 155460 3392
rect 156604 3340 156656 3392
rect 160100 3340 160152 3392
rect 161296 3340 161348 3392
rect 181444 3340 181496 3392
rect 215300 3340 215352 3392
rect 222752 3340 222804 3392
rect 233332 3340 233384 3392
rect 324320 3340 324372 3392
rect 144736 3272 144788 3324
rect 148324 3272 148376 3324
rect 188528 3272 188580 3324
rect 218152 3272 218204 3324
rect 225144 3272 225196 3324
rect 234804 3272 234856 3324
rect 248512 3272 248564 3324
rect 257068 3272 257120 3324
rect 321560 3272 321612 3324
rect 422576 3272 422628 3324
rect 423772 3340 423824 3392
rect 424968 3340 425020 3392
rect 431960 3340 432012 3392
rect 433248 3340 433300 3392
rect 440332 3340 440384 3392
rect 441528 3340 441580 3392
rect 429660 3272 429712 3324
rect 473360 3476 473412 3528
rect 474188 3476 474240 3528
rect 489920 3476 489972 3528
rect 490748 3476 490800 3528
rect 498200 3476 498252 3528
rect 499028 3476 499080 3528
rect 514760 3476 514812 3528
rect 515588 3476 515640 3528
rect 523040 3476 523092 3528
rect 523868 3476 523920 3528
rect 539600 3476 539652 3528
rect 540428 3476 540480 3528
rect 564440 3476 564492 3528
rect 565268 3476 565320 3528
rect 570604 3476 570656 3528
rect 571524 3476 571576 3528
rect 479340 3340 479392 3392
rect 581000 3408 581052 3460
rect 192024 3204 192076 3256
rect 219716 3204 219768 3256
rect 226340 3204 226392 3256
rect 236000 3204 236052 3256
rect 317512 3204 317564 3256
rect 415400 3204 415452 3256
rect 415492 3204 415544 3256
rect 416688 3204 416740 3256
rect 151820 3136 151872 3188
rect 155224 3136 155276 3188
rect 221556 3136 221608 3188
rect 233608 3136 233660 3188
rect 390560 3136 390612 3188
rect 392032 3136 392084 3188
rect 398932 3136 398984 3188
rect 400128 3136 400180 3188
rect 407212 3136 407264 3188
rect 408408 3136 408460 3188
rect 205088 3068 205140 3120
rect 226524 3068 226576 3120
rect 137652 3000 137704 3052
rect 140044 3000 140096 3052
rect 234620 3000 234672 3052
rect 238944 3000 238996 3052
rect 248604 3000 248656 3052
rect 255872 3000 255924 3052
rect 571984 3000 572036 3052
rect 573916 3000 573968 3052
rect 148324 2932 148376 2984
rect 152464 2932 152516 2984
rect 233424 2864 233476 2916
rect 238024 2864 238076 2916
rect 448520 1912 448572 1964
rect 449808 1912 449860 1964
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3330 606112 3386 606121
rect 3330 606047 3386 606056
rect 3344 605878 3372 606047
rect 3332 605872 3384 605878
rect 3332 605814 3384 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 2870 475688 2926 475697
rect 2870 475623 2926 475632
rect 2884 474774 2912 475623
rect 2872 474768 2924 474774
rect 2872 474710 2924 474716
rect 2778 423600 2834 423609
rect 2778 423535 2780 423544
rect 2832 423535 2834 423544
rect 2780 423506 2832 423512
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3344 409902 3372 410479
rect 3332 409896 3384 409902
rect 3332 409838 3384 409844
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 3436 362302 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 362370 3556 619103
rect 3606 566944 3662 566953
rect 3606 566879 3662 566888
rect 3620 362506 3648 566879
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3712 362574 3740 553823
rect 3790 501800 3846 501809
rect 3790 501735 3846 501744
rect 3804 362642 3832 501735
rect 3882 462632 3938 462641
rect 3882 462567 3938 462576
rect 3896 362710 3924 462567
rect 3974 449576 4030 449585
rect 3974 449511 4030 449520
rect 3988 362778 4016 449511
rect 4804 423564 4856 423570
rect 4804 423506 4856 423512
rect 4066 397488 4122 397497
rect 4066 397423 4122 397432
rect 4080 362846 4108 397423
rect 4816 367810 4844 423506
rect 4804 367804 4856 367810
rect 4804 367746 4856 367752
rect 4068 362840 4120 362846
rect 4068 362782 4120 362788
rect 3976 362772 4028 362778
rect 3976 362714 4028 362720
rect 3884 362704 3936 362710
rect 3884 362646 3936 362652
rect 3792 362636 3844 362642
rect 3792 362578 3844 362584
rect 3700 362568 3752 362574
rect 3700 362510 3752 362516
rect 3608 362500 3660 362506
rect 3608 362442 3660 362448
rect 3516 362364 3568 362370
rect 3516 362306 3568 362312
rect 3424 362296 3476 362302
rect 3424 362238 3476 362244
rect 6932 362234 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 13820 371272 13872 371278
rect 13820 371214 13872 371220
rect 13832 369170 13860 371214
rect 13820 369164 13872 369170
rect 13820 369106 13872 369112
rect 23492 362438 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 40052 366382 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 40040 366376 40092 366382
rect 40040 366318 40092 366324
rect 71792 362914 71820 702986
rect 89180 702434 89208 703520
rect 88352 702406 89208 702434
rect 71780 362908 71832 362914
rect 71780 362850 71832 362856
rect 23480 362432 23532 362438
rect 23480 362374 23532 362380
rect 6920 362228 6972 362234
rect 6920 362170 6972 362176
rect 88352 362166 88380 702406
rect 93124 683188 93176 683194
rect 93124 683130 93176 683136
rect 93136 370530 93164 683130
rect 93124 370524 93176 370530
rect 93124 370466 93176 370472
rect 104912 365022 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 136652 371890 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702434 154160 703520
rect 153212 702406 154160 702434
rect 136640 371884 136692 371890
rect 136640 371826 136692 371832
rect 104900 365016 104952 365022
rect 104900 364958 104952 364964
rect 88340 362160 88392 362166
rect 88340 362102 88392 362108
rect 153212 362098 153240 702406
rect 170324 700330 170352 703520
rect 202800 700330 202828 703520
rect 170312 700324 170364 700330
rect 170312 700266 170364 700272
rect 192484 700324 192536 700330
rect 192484 700266 192536 700272
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 192496 363662 192524 700266
rect 211160 409896 211212 409902
rect 211160 409838 211212 409844
rect 205640 369164 205692 369170
rect 205640 369106 205692 369112
rect 192484 363656 192536 363662
rect 192484 363598 192536 363604
rect 153200 362092 153252 362098
rect 153200 362034 153252 362040
rect 186964 360528 187016 360534
rect 186964 360470 187016 360476
rect 195704 360528 195756 360534
rect 195704 360470 195756 360476
rect 4804 360460 4856 360466
rect 4804 360402 4856 360408
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 3424 343664 3476 343670
rect 3424 343606 3476 343612
rect 2780 319864 2832 319870
rect 2780 319806 2832 319812
rect 2792 319297 2820 319806
rect 2778 319288 2834 319297
rect 2778 319223 2834 319232
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 3068 293185 3096 293898
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 3436 254153 3464 343606
rect 4816 319870 4844 360402
rect 7564 334008 7616 334014
rect 7564 333950 7616 333956
rect 4804 319864 4856 319870
rect 4804 319806 4856 319812
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 4804 303680 4856 303686
rect 4804 303622 4856 303628
rect 3516 267708 3568 267714
rect 3516 267650 3568 267656
rect 3528 267209 3556 267650
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3608 253972 3660 253978
rect 3608 253914 3660 253920
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3516 225004 3568 225010
rect 3516 224946 3568 224952
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3424 194608 3476 194614
rect 3424 194550 3476 194556
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 164212 3384 164218
rect 3332 164154 3384 164160
rect 3344 162897 3372 164154
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3344 149841 3372 150350
rect 3330 149832 3386 149841
rect 3330 149767 3386 149776
rect 3056 137964 3108 137970
rect 3056 137906 3108 137912
rect 3068 136785 3096 137906
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 3332 110900 3384 110906
rect 3332 110842 3384 110848
rect 3344 110673 3372 110842
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3436 19417 3464 194550
rect 3528 58585 3556 224946
rect 3620 97617 3648 253914
rect 4816 215286 4844 303622
rect 7576 267714 7604 333950
rect 22744 324352 22796 324358
rect 22744 324294 22796 324300
rect 14464 274712 14516 274718
rect 14464 274654 14516 274660
rect 7564 267708 7616 267714
rect 7564 267650 7616 267656
rect 7564 244316 7616 244322
rect 7564 244258 7616 244264
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 7576 110906 7604 244258
rect 14476 164218 14504 274654
rect 21364 213988 21416 213994
rect 21364 213930 21416 213936
rect 14464 164212 14516 164218
rect 14464 164154 14516 164160
rect 7564 110900 7616 110906
rect 7564 110842 7616 110848
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 21376 71738 21404 213930
rect 22756 189038 22784 324294
rect 186976 306338 187004 360470
rect 191104 360392 191156 360398
rect 191104 360334 191156 360340
rect 188344 360256 188396 360262
rect 188344 360198 188396 360204
rect 186964 306332 187016 306338
rect 186964 306274 187016 306280
rect 188356 293962 188384 360198
rect 189722 354784 189778 354793
rect 189722 354719 189778 354728
rect 189078 344312 189134 344321
rect 189078 344247 189134 344256
rect 189092 343670 189120 344247
rect 189080 343664 189132 343670
rect 189080 343606 189132 343612
rect 189078 334384 189134 334393
rect 189078 334319 189134 334328
rect 189092 334014 189120 334319
rect 189080 334008 189132 334014
rect 189080 333950 189132 333956
rect 189078 324456 189134 324465
rect 189078 324391 189134 324400
rect 189092 324358 189120 324391
rect 189080 324352 189132 324358
rect 189080 324294 189132 324300
rect 189078 304328 189134 304337
rect 189078 304263 189134 304272
rect 189092 303686 189120 304263
rect 189080 303680 189132 303686
rect 189080 303622 189132 303628
rect 188344 293956 188396 293962
rect 188344 293898 188396 293904
rect 189078 274816 189134 274825
rect 189078 274751 189134 274760
rect 189092 274718 189120 274751
rect 189080 274712 189132 274718
rect 189080 274654 189132 274660
rect 189078 254280 189134 254289
rect 189078 254215 189134 254224
rect 189092 253978 189120 254215
rect 189080 253972 189132 253978
rect 189080 253914 189132 253920
rect 189078 244352 189134 244361
rect 189078 244287 189080 244296
rect 189132 244287 189134 244296
rect 189080 244258 189132 244264
rect 189736 241466 189764 354719
rect 191116 346390 191144 360334
rect 191748 360324 191800 360330
rect 191748 360266 191800 360272
rect 191760 358766 191788 360266
rect 193220 360256 193272 360262
rect 193220 360198 193272 360204
rect 193232 359924 193260 360198
rect 195716 359924 195744 360470
rect 198280 360460 198332 360466
rect 198280 360402 198332 360408
rect 198292 359924 198320 360402
rect 200856 360392 200908 360398
rect 200856 360334 200908 360340
rect 200868 359924 200896 360334
rect 203432 360324 203484 360330
rect 203432 360266 203484 360272
rect 203444 359924 203472 360266
rect 205652 359938 205680 369106
rect 208584 362840 208636 362846
rect 208584 362782 208636 362788
rect 205652 359910 206034 359938
rect 208596 359924 208624 362782
rect 211172 359924 211200 409838
rect 213184 367804 213236 367810
rect 213184 367746 213236 367752
rect 213196 359938 213224 367746
rect 218072 362846 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 235184 700330 235212 703520
rect 220084 700324 220136 700330
rect 220084 700266 220136 700272
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 220096 476814 220124 700266
rect 267660 697610 267688 703520
rect 282184 700324 282236 700330
rect 282184 700266 282236 700272
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 246304 656940 246356 656946
rect 246304 656882 246356 656888
rect 244280 632120 244332 632126
rect 244280 632062 244332 632068
rect 238024 605872 238076 605878
rect 238024 605814 238076 605820
rect 235264 579692 235316 579698
rect 235264 579634 235316 579640
rect 228364 527196 228416 527202
rect 228364 527138 228416 527144
rect 226340 514820 226392 514826
rect 226340 514762 226392 514768
rect 220084 476808 220136 476814
rect 220084 476750 220136 476756
rect 220084 474768 220136 474774
rect 220084 474710 220136 474716
rect 220096 362982 220124 474710
rect 220084 362976 220136 362982
rect 220084 362918 220136 362924
rect 221372 362976 221424 362982
rect 221372 362918 221424 362924
rect 218060 362840 218112 362846
rect 218060 362782 218112 362788
rect 216220 362772 216272 362778
rect 216220 362714 216272 362720
rect 213196 359910 213670 359938
rect 216232 359924 216260 362714
rect 218796 362704 218848 362710
rect 218796 362646 218848 362652
rect 218808 359924 218836 362646
rect 221384 359924 221412 362918
rect 223948 362636 224000 362642
rect 223948 362578 224000 362584
rect 223960 359924 223988 362578
rect 226352 359938 226380 514762
rect 228376 363254 228404 527138
rect 228364 363248 228416 363254
rect 228364 363190 228416 363196
rect 229100 363248 229152 363254
rect 229100 363190 229152 363196
rect 226352 359910 226550 359938
rect 229112 359924 229140 363190
rect 235276 362982 235304 579634
rect 238036 363254 238064 605814
rect 238024 363248 238076 363254
rect 238024 363190 238076 363196
rect 239312 363248 239364 363254
rect 239312 363190 239364 363196
rect 235264 362976 235316 362982
rect 235264 362918 235316 362924
rect 236736 362976 236788 362982
rect 236736 362918 236788 362924
rect 231676 362568 231728 362574
rect 231676 362510 231728 362516
rect 231688 359924 231716 362510
rect 234160 362500 234212 362506
rect 234160 362442 234212 362448
rect 234172 359924 234200 362442
rect 236748 359924 236776 362918
rect 239324 359924 239352 363190
rect 241888 362364 241940 362370
rect 241888 362306 241940 362312
rect 241900 359924 241928 362306
rect 244292 359938 244320 632062
rect 246316 362982 246344 656882
rect 251824 370524 251876 370530
rect 251824 370466 251876 370472
rect 246304 362976 246356 362982
rect 246304 362918 246356 362924
rect 247040 362976 247092 362982
rect 247040 362918 247092 362924
rect 244292 359910 244490 359938
rect 247052 359924 247080 362918
rect 249616 362296 249668 362302
rect 249616 362238 249668 362244
rect 249628 359924 249656 362238
rect 251836 359938 251864 370466
rect 259828 366376 259880 366382
rect 259828 366318 259880 366324
rect 257252 362432 257304 362438
rect 257252 362374 257304 362380
rect 254676 362228 254728 362234
rect 254676 362170 254728 362176
rect 251836 359910 252218 359938
rect 254688 359924 254716 362170
rect 257264 359924 257292 362374
rect 259840 359924 259868 366318
rect 262404 362908 262456 362914
rect 262404 362850 262456 362856
rect 262416 359924 262444 362850
rect 266372 362234 266400 697546
rect 277400 476808 277452 476814
rect 277400 476750 277452 476756
rect 269672 371884 269724 371890
rect 269672 371826 269724 371832
rect 267556 365016 267608 365022
rect 267556 364958 267608 364964
rect 266360 362228 266412 362234
rect 266360 362170 266412 362176
rect 264980 362160 265032 362166
rect 264980 362102 265032 362108
rect 264992 359924 265020 362102
rect 267568 359924 267596 364958
rect 269684 359938 269712 371826
rect 275192 363656 275244 363662
rect 275192 363598 275244 363604
rect 272708 362092 272760 362098
rect 272708 362034 272760 362040
rect 269684 359910 270158 359938
rect 272720 359924 272748 362034
rect 275204 359924 275232 363598
rect 277412 359938 277440 476750
rect 280344 362840 280396 362846
rect 280344 362782 280396 362788
rect 277412 359910 277794 359938
rect 280356 359924 280384 362782
rect 282196 361894 282224 700266
rect 283852 700126 283880 703520
rect 292580 700936 292632 700942
rect 292580 700878 292632 700884
rect 291844 700324 291896 700330
rect 291844 700266 291896 700272
rect 283840 700120 283892 700126
rect 283840 700062 283892 700068
rect 284944 700120 284996 700126
rect 284944 700062 284996 700068
rect 284956 362914 284984 700062
rect 284944 362908 284996 362914
rect 284944 362850 284996 362856
rect 288072 362908 288124 362914
rect 288072 362850 288124 362856
rect 285496 362228 285548 362234
rect 285496 362170 285548 362176
rect 282184 361888 282236 361894
rect 282184 361830 282236 361836
rect 282920 361888 282972 361894
rect 282920 361830 282972 361836
rect 282932 359924 282960 361830
rect 285508 359924 285536 362170
rect 288084 359924 288112 362850
rect 291856 361894 291884 700266
rect 292592 383654 292620 700878
rect 295340 700868 295392 700874
rect 295340 700810 295392 700816
rect 292592 383626 292896 383654
rect 290648 361888 290700 361894
rect 290648 361830 290700 361836
rect 291844 361888 291896 361894
rect 291844 361830 291896 361836
rect 290660 359924 290688 361830
rect 292868 359938 292896 383626
rect 295352 359938 295380 700810
rect 298100 700800 298152 700806
rect 298100 700742 298152 700748
rect 298112 359938 298140 700742
rect 300136 700330 300164 703520
rect 332520 700942 332548 703520
rect 332508 700936 332560 700942
rect 332508 700878 332560 700884
rect 348804 700874 348832 703520
rect 348792 700868 348844 700874
rect 348792 700810 348844 700816
rect 364996 700806 365024 703520
rect 364984 700800 365036 700806
rect 364984 700742 365036 700748
rect 397472 700738 397500 703520
rect 300860 700732 300912 700738
rect 300860 700674 300912 700680
rect 397460 700732 397512 700738
rect 397460 700674 397512 700680
rect 300124 700324 300176 700330
rect 300124 700266 300176 700272
rect 292868 359910 293250 359938
rect 295352 359910 295734 359938
rect 298112 359910 298310 359938
rect 300872 359924 300900 700674
rect 413664 700670 413692 703520
rect 302240 700664 302292 700670
rect 302240 700606 302292 700612
rect 413652 700664 413704 700670
rect 413652 700606 413704 700612
rect 302252 383654 302280 700606
rect 429856 700602 429884 703520
rect 305000 700596 305052 700602
rect 305000 700538 305052 700544
rect 429844 700596 429896 700602
rect 429844 700538 429896 700544
rect 305012 383654 305040 700538
rect 462332 700534 462360 703520
rect 307760 700528 307812 700534
rect 307760 700470 307812 700476
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 307772 383654 307800 700470
rect 478524 700466 478552 703520
rect 310520 700460 310572 700466
rect 310520 700402 310572 700408
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 310532 383654 310560 700402
rect 316040 700392 316092 700398
rect 316040 700334 316092 700340
rect 302252 383626 303016 383654
rect 305012 383626 305592 383654
rect 307772 383626 308168 383654
rect 310532 383626 310744 383654
rect 302988 359938 303016 383626
rect 305564 359938 305592 383626
rect 308140 359938 308168 383626
rect 310716 359938 310744 383626
rect 313648 362296 313700 362302
rect 313648 362238 313700 362244
rect 302988 359910 303462 359938
rect 305564 359910 306038 359938
rect 308140 359910 308614 359938
rect 310716 359910 311190 359938
rect 313660 359924 313688 362238
rect 316052 359938 316080 700334
rect 318800 700324 318852 700330
rect 318800 700266 318852 700272
rect 316052 359910 316250 359938
rect 318812 359924 318840 700266
rect 322940 696992 322992 696998
rect 322940 696934 322992 696940
rect 322952 383654 322980 696934
rect 325700 683188 325752 683194
rect 325700 683130 325752 683136
rect 325712 383654 325740 683130
rect 328460 670744 328512 670750
rect 328460 670686 328512 670692
rect 328472 383654 328500 670686
rect 331220 643136 331272 643142
rect 331220 643078 331272 643084
rect 331232 383654 331260 643078
rect 333980 630692 334032 630698
rect 333980 630634 334032 630640
rect 322952 383626 323624 383654
rect 325712 383626 326200 383654
rect 328472 383626 328776 383654
rect 331232 383626 331352 383654
rect 321376 362228 321428 362234
rect 321376 362170 321428 362176
rect 321388 359924 321416 362170
rect 323596 359938 323624 383626
rect 326172 359938 326200 383626
rect 328748 359938 328776 383626
rect 331324 359938 331352 383626
rect 333992 359938 334020 630634
rect 336740 616888 336792 616894
rect 336740 616830 336792 616836
rect 323596 359910 323978 359938
rect 326172 359910 326554 359938
rect 328748 359910 329130 359938
rect 331324 359910 331706 359938
rect 333992 359910 334190 359938
rect 336752 359924 336780 616830
rect 338120 590708 338172 590714
rect 338120 590650 338172 590656
rect 338132 383654 338160 590650
rect 340880 576904 340932 576910
rect 340880 576846 340932 576852
rect 340892 383654 340920 576846
rect 343640 563100 343692 563106
rect 343640 563042 343692 563048
rect 343652 383654 343680 563042
rect 346400 536852 346452 536858
rect 346400 536794 346452 536800
rect 346412 383654 346440 536794
rect 349160 524476 349212 524482
rect 349160 524418 349212 524424
rect 338132 383626 338896 383654
rect 340892 383626 341472 383654
rect 343652 383626 344048 383654
rect 346412 383626 346624 383654
rect 338868 359938 338896 383626
rect 341444 359938 341472 383626
rect 344020 359938 344048 383626
rect 346596 359938 346624 383626
rect 349172 359938 349200 524418
rect 351920 510672 351972 510678
rect 351920 510614 351972 510620
rect 351932 359938 351960 510614
rect 354680 484424 354732 484430
rect 354680 484366 354732 484372
rect 338868 359910 339342 359938
rect 341444 359910 341918 359938
rect 344020 359910 344494 359938
rect 346596 359910 347070 359938
rect 349172 359910 349646 359938
rect 351932 359910 352222 359938
rect 354692 359924 354720 484366
rect 356060 470620 356112 470626
rect 356060 470562 356112 470568
rect 356072 383654 356100 470562
rect 358820 456816 358872 456822
rect 358820 456758 358872 456764
rect 358832 383654 358860 456758
rect 361580 430636 361632 430642
rect 361580 430578 361632 430584
rect 361592 383654 361620 430578
rect 364340 418192 364392 418198
rect 364340 418134 364392 418140
rect 364352 383654 364380 418134
rect 367100 404388 367152 404394
rect 367100 404330 367152 404336
rect 367112 383654 367140 404330
rect 356072 383626 356928 383654
rect 358832 383626 359504 383654
rect 361592 383626 362080 383654
rect 364352 383626 364656 383654
rect 367112 383626 367232 383654
rect 356900 359938 356928 383626
rect 359476 359938 359504 383626
rect 362052 359938 362080 383626
rect 364628 359938 364656 383626
rect 367204 359938 367232 383626
rect 369860 378208 369912 378214
rect 369860 378150 369912 378156
rect 369872 359938 369900 378150
rect 372712 364404 372764 364410
rect 372712 364346 372764 364352
rect 356900 359910 357282 359938
rect 359476 359910 359858 359938
rect 362052 359910 362434 359938
rect 364628 359910 365010 359938
rect 367204 359910 367586 359938
rect 369872 359910 370162 359938
rect 372724 359924 372752 364346
rect 494072 362302 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 494060 362296 494112 362302
rect 494060 362238 494112 362244
rect 558932 362234 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 558920 362228 558972 362234
rect 558920 362170 558972 362176
rect 382924 361956 382976 361962
rect 382924 361898 382976 361904
rect 479524 361956 479576 361962
rect 479524 361898 479576 361904
rect 377772 361752 377824 361758
rect 377772 361694 377824 361700
rect 375196 361684 375248 361690
rect 375196 361626 375248 361632
rect 375208 359924 375236 361626
rect 377784 359924 377812 361694
rect 380348 361616 380400 361622
rect 380348 361558 380400 361564
rect 380360 359924 380388 361558
rect 382936 359924 382964 361898
rect 388076 361888 388128 361894
rect 388076 361830 388128 361836
rect 385500 361820 385552 361826
rect 385500 361762 385552 361768
rect 385512 359924 385540 361762
rect 388088 359924 388116 361830
rect 390928 359440 390980 359446
rect 390678 359388 390928 359394
rect 390678 359382 390980 359388
rect 391848 359440 391900 359446
rect 391848 359382 391900 359388
rect 390678 359366 390968 359382
rect 391860 358834 391888 359382
rect 391848 358828 391900 358834
rect 391848 358770 391900 358776
rect 406384 358828 406436 358834
rect 406384 358770 406436 358776
rect 191748 358760 191800 358766
rect 191748 358702 191800 358708
rect 394146 354784 394202 354793
rect 394146 354719 394202 354728
rect 191104 346384 191156 346390
rect 191104 346326 191156 346332
rect 394054 344312 394110 344321
rect 394054 344247 394110 344256
rect 393962 334384 394018 334393
rect 393962 334319 394018 334328
rect 190090 314800 190146 314809
rect 190090 314735 190146 314744
rect 189998 294400 190054 294409
rect 189998 294335 190054 294344
rect 189906 264344 189962 264353
rect 189906 264279 189962 264288
rect 189724 241460 189776 241466
rect 189724 241402 189776 241408
rect 189814 234696 189870 234705
rect 189814 234631 189870 234640
rect 189078 225040 189134 225049
rect 189078 224975 189080 224984
rect 189132 224975 189134 224984
rect 189080 224946 189132 224952
rect 189078 214296 189134 214305
rect 189078 214231 189134 214240
rect 189092 213994 189120 214231
rect 189080 213988 189132 213994
rect 189080 213930 189132 213936
rect 189722 204368 189778 204377
rect 189722 204303 189778 204312
rect 189078 194712 189134 194721
rect 189078 194647 189134 194656
rect 189092 194614 189120 194647
rect 189080 194608 189132 194614
rect 189080 194550 189132 194556
rect 22744 189032 22796 189038
rect 22744 188974 22796 188980
rect 188344 177676 188396 177682
rect 188344 177618 188396 177624
rect 184940 177540 184992 177546
rect 184940 177482 184992 177488
rect 176660 177472 176712 177478
rect 176660 177414 176712 177420
rect 141424 177404 141476 177410
rect 141424 177346 141476 177352
rect 134524 177336 134576 177342
rect 134524 177278 134576 177284
rect 125600 175976 125652 175982
rect 125600 175918 125652 175924
rect 21364 71732 21416 71738
rect 21364 71674 21416 71680
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125612 354 125640 175918
rect 129740 156664 129792 156670
rect 129740 156606 129792 156612
rect 129752 16574 129780 156606
rect 129752 16546 130608 16574
rect 129004 10328 129056 10334
rect 129004 10270 129056 10276
rect 128176 4072 128228 4078
rect 128176 4014 128228 4020
rect 126980 3528 127032 3534
rect 126980 3470 127032 3476
rect 126992 480 127020 3470
rect 128188 480 128216 4014
rect 129016 3534 129044 10270
rect 129372 4820 129424 4826
rect 129372 4762 129424 4768
rect 129004 3528 129056 3534
rect 129004 3470 129056 3476
rect 129384 480 129412 4762
rect 130580 480 130608 16546
rect 132960 4888 133012 4894
rect 132960 4830 133012 4836
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 131776 480 131804 3402
rect 132972 480 133000 4830
rect 134536 4078 134564 177278
rect 137284 155236 137336 155242
rect 137284 155178 137336 155184
rect 136456 4956 136508 4962
rect 136456 4898 136508 4904
rect 134524 4072 134576 4078
rect 134524 4014 134576 4020
rect 134156 3528 134208 3534
rect 134156 3470 134208 3476
rect 134168 480 134196 3470
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 135272 480 135300 3334
rect 136468 480 136496 4898
rect 137296 3534 137324 155178
rect 140044 153876 140096 153882
rect 140044 153818 140096 153824
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 138846 3360 138902 3369
rect 138846 3295 138902 3304
rect 137652 3052 137704 3058
rect 137652 2994 137704 3000
rect 137664 480 137692 2994
rect 138860 480 138888 3295
rect 140056 3058 140084 153818
rect 140136 5024 140188 5030
rect 140136 4966 140188 4972
rect 140044 3052 140096 3058
rect 140044 2994 140096 3000
rect 140148 2530 140176 4966
rect 141240 4140 141292 4146
rect 141240 4082 141292 4088
rect 140056 2502 140176 2530
rect 140056 480 140084 2502
rect 141252 480 141280 4082
rect 141436 3398 141464 177346
rect 160100 174616 160152 174622
rect 160100 174558 160152 174564
rect 155224 174548 155276 174554
rect 155224 174490 155276 174496
rect 142804 171828 142856 171834
rect 142804 171770 142856 171776
rect 142816 4146 142844 171770
rect 143540 170400 143592 170406
rect 143540 170342 143592 170348
rect 142804 4140 142856 4146
rect 142804 4082 142856 4088
rect 142436 3528 142488 3534
rect 142436 3470 142488 3476
rect 141424 3392 141476 3398
rect 141424 3334 141476 3340
rect 142448 480 142476 3470
rect 143552 480 143580 170342
rect 146300 169040 146352 169046
rect 146300 168982 146352 168988
rect 146312 16574 146340 168982
rect 150440 167680 150492 167686
rect 150440 167622 150492 167628
rect 148324 152516 148376 152522
rect 148324 152458 148376 152464
rect 146312 16546 147168 16574
rect 145932 3596 145984 3602
rect 145932 3538 145984 3544
rect 144736 3324 144788 3330
rect 144736 3266 144788 3272
rect 144748 480 144776 3266
rect 145944 480 145972 3538
rect 147140 480 147168 16546
rect 148336 3330 148364 152458
rect 150452 16574 150480 167622
rect 152464 151088 152516 151094
rect 152464 151030 152516 151036
rect 150452 16546 150664 16574
rect 149520 3664 149572 3670
rect 149520 3606 149572 3612
rect 148324 3324 148376 3330
rect 148324 3266 148376 3272
rect 148324 2984 148376 2990
rect 148324 2926 148376 2932
rect 148336 480 148364 2926
rect 149532 480 149560 3606
rect 150636 480 150664 16546
rect 151820 3188 151872 3194
rect 151820 3130 151872 3136
rect 151832 480 151860 3130
rect 152476 2990 152504 151030
rect 154212 8968 154264 8974
rect 154212 8910 154264 8916
rect 153016 3732 153068 3738
rect 153016 3674 153068 3680
rect 152464 2984 152516 2990
rect 152464 2926 152516 2932
rect 153028 480 153056 3674
rect 154224 480 154252 8910
rect 155236 3194 155264 174490
rect 158720 173188 158772 173194
rect 158720 173130 158772 173136
rect 157340 166320 157392 166326
rect 157340 166262 157392 166268
rect 156604 148368 156656 148374
rect 156604 148310 156656 148316
rect 156616 3398 156644 148310
rect 157352 16574 157380 166262
rect 158732 16574 158760 173130
rect 157352 16546 157840 16574
rect 158732 16546 158944 16574
rect 156696 3800 156748 3806
rect 156696 3742 156748 3748
rect 155408 3392 155460 3398
rect 155408 3334 155460 3340
rect 156604 3392 156656 3398
rect 156604 3334 156656 3340
rect 155224 3188 155276 3194
rect 155224 3130 155276 3136
rect 155420 480 155448 3334
rect 156708 1986 156736 3742
rect 156616 1958 156736 1986
rect 156616 480 156644 1958
rect 157812 480 157840 16546
rect 158916 480 158944 16546
rect 160112 3398 160140 174558
rect 164240 173256 164292 173262
rect 164240 173198 164292 173204
rect 161480 164892 161532 164898
rect 161480 164834 161532 164840
rect 161492 16574 161520 164834
rect 164252 16574 164280 173198
rect 168380 171896 168432 171902
rect 168380 171838 168432 171844
rect 165620 163532 165672 163538
rect 165620 163474 165672 163480
rect 165632 16574 165660 163474
rect 161492 16546 162072 16574
rect 164252 16546 164464 16574
rect 165632 16546 166120 16574
rect 160192 3868 160244 3874
rect 160192 3810 160244 3816
rect 160100 3392 160152 3398
rect 160100 3334 160152 3340
rect 160204 1986 160232 3810
rect 161296 3392 161348 3398
rect 161296 3334 161348 3340
rect 160112 1958 160232 1986
rect 160112 480 160140 1958
rect 161308 480 161336 3334
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162044 354 162072 16546
rect 163688 3936 163740 3942
rect 163688 3878 163740 3884
rect 163700 480 163728 3878
rect 162462 354 162574 480
rect 162044 326 162574 354
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164436 354 164464 16546
rect 166092 480 166120 16546
rect 167184 4072 167236 4078
rect 167184 4014 167236 4020
rect 167196 480 167224 4014
rect 168392 480 168420 171838
rect 172520 162172 172572 162178
rect 172520 162114 172572 162120
rect 172532 16574 172560 162114
rect 172532 16546 172744 16574
rect 169576 11756 169628 11762
rect 169576 11698 169628 11704
rect 169588 480 169616 11698
rect 171968 7608 172020 7614
rect 171968 7550 172020 7556
rect 170772 4004 170824 4010
rect 170772 3946 170824 3952
rect 170784 480 170812 3946
rect 171980 480 172008 7550
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 172716 354 172744 16546
rect 176672 11830 176700 177414
rect 176752 160744 176804 160750
rect 176752 160686 176804 160692
rect 176660 11824 176712 11830
rect 176660 11766 176712 11772
rect 176764 6914 176792 160686
rect 179420 159384 179472 159390
rect 179420 159326 179472 159332
rect 179432 16574 179460 159326
rect 183560 158024 183612 158030
rect 183560 157966 183612 157972
rect 183572 16574 183600 157966
rect 179432 16546 180288 16574
rect 183572 16546 183784 16574
rect 177856 11824 177908 11830
rect 177856 11766 177908 11772
rect 176672 6886 176792 6914
rect 175464 5092 175516 5098
rect 175464 5034 175516 5040
rect 174268 4140 174320 4146
rect 174268 4082 174320 4088
rect 174280 480 174308 4082
rect 175476 480 175504 5034
rect 176672 480 176700 6886
rect 177868 480 177896 11766
rect 179052 5160 179104 5166
rect 179052 5102 179104 5108
rect 179064 480 179092 5102
rect 180260 480 180288 16546
rect 182548 5228 182600 5234
rect 182548 5170 182600 5176
rect 181444 3392 181496 3398
rect 181444 3334 181496 3340
rect 181456 480 181484 3334
rect 182560 480 182588 5170
rect 183756 480 183784 16546
rect 184952 480 184980 177482
rect 186320 170468 186372 170474
rect 186320 170410 186372 170416
rect 186332 16574 186360 170410
rect 186332 16546 186912 16574
rect 186136 6180 186188 6186
rect 186136 6122 186188 6128
rect 186148 480 186176 6122
rect 173134 354 173246 480
rect 172716 326 173246 354
rect 173134 -960 173246 326
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 186884 354 186912 16546
rect 188356 8974 188384 177618
rect 188344 8968 188396 8974
rect 188344 8910 188396 8916
rect 189736 6866 189764 204303
rect 189828 45558 189856 234631
rect 189920 85542 189948 264279
rect 190012 137970 190040 294335
rect 190104 202842 190132 314735
rect 190182 284336 190238 284345
rect 190182 284271 190238 284280
rect 190092 202836 190144 202842
rect 190092 202778 190144 202784
rect 190090 185056 190146 185065
rect 190090 184991 190146 185000
rect 190000 137964 190052 137970
rect 190000 137906 190052 137912
rect 189908 85536 189960 85542
rect 189908 85478 189960 85484
rect 189816 45552 189868 45558
rect 189816 45494 189868 45500
rect 190104 33114 190132 184991
rect 190196 150414 190224 284271
rect 393778 244624 393834 244633
rect 393778 244559 393780 244568
rect 393832 244559 393834 244568
rect 393780 244530 393832 244536
rect 393976 206990 394004 334319
rect 394068 219434 394096 344247
rect 394160 233238 394188 354719
rect 394606 324456 394662 324465
rect 394606 324391 394662 324400
rect 394330 314800 394386 314809
rect 394330 314735 394332 314744
rect 394384 314735 394386 314744
rect 394332 314706 394384 314712
rect 394330 304328 394386 304337
rect 394330 304263 394386 304272
rect 394344 303686 394372 304263
rect 394332 303680 394384 303686
rect 394332 303622 394384 303628
rect 394514 294400 394570 294409
rect 394514 294335 394570 294344
rect 394422 284608 394478 284617
rect 394422 284543 394424 284552
rect 394476 284543 394478 284552
rect 394424 284514 394476 284520
rect 394422 274816 394478 274825
rect 394422 274751 394478 274760
rect 394436 274718 394464 274751
rect 394424 274712 394476 274718
rect 394424 274654 394476 274660
rect 394422 264344 394478 264353
rect 394422 264279 394478 264288
rect 394330 254280 394386 254289
rect 394330 254215 394386 254224
rect 394238 234696 394294 234705
rect 394238 234631 394294 234640
rect 394148 233232 394200 233238
rect 394148 233174 394200 233180
rect 394146 225040 394202 225049
rect 394146 224975 394202 224984
rect 394056 219428 394108 219434
rect 394056 219370 394108 219376
rect 394054 214432 394110 214441
rect 394054 214367 394110 214376
rect 394068 213994 394096 214367
rect 394056 213988 394108 213994
rect 394056 213930 394108 213936
rect 393964 206984 394016 206990
rect 393964 206926 394016 206932
rect 394054 204368 394110 204377
rect 394054 204303 394110 204312
rect 393962 194712 394018 194721
rect 393962 194647 394018 194656
rect 356086 180254 356376 180282
rect 382398 180254 382596 180282
rect 191944 180118 192234 180146
rect 192312 180118 192694 180146
rect 193246 180118 193352 180146
rect 191104 177608 191156 177614
rect 191104 177550 191156 177556
rect 190460 169108 190512 169114
rect 190460 169050 190512 169056
rect 190184 150408 190236 150414
rect 190184 150350 190236 150356
rect 190092 33108 190144 33114
rect 190092 33050 190144 33056
rect 189724 6860 189776 6866
rect 189724 6802 189776 6808
rect 189724 5296 189776 5302
rect 189724 5238 189776 5244
rect 188528 3324 188580 3330
rect 188528 3266 188580 3272
rect 188540 480 188568 3266
rect 189736 480 189764 5238
rect 187302 354 187414 480
rect 186884 326 187414 354
rect 187302 -960 187414 326
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190472 354 190500 169050
rect 191116 7614 191144 177550
rect 191944 10334 191972 180118
rect 192312 177342 192340 180118
rect 192300 177336 192352 177342
rect 192300 177278 192352 177284
rect 192484 176724 192536 176730
rect 192484 176666 192536 176672
rect 192496 156670 192524 176666
rect 192484 156664 192536 156670
rect 192484 156606 192536 156612
rect 191932 10328 191984 10334
rect 191932 10270 191984 10276
rect 191104 7608 191156 7614
rect 191104 7550 191156 7556
rect 193324 4826 193352 180118
rect 193416 180118 193706 180146
rect 193876 180118 194258 180146
rect 194612 180118 194810 180146
rect 194888 180118 195270 180146
rect 195440 180118 195822 180146
rect 195992 180118 196282 180146
rect 196452 180118 196834 180146
rect 197386 180118 197492 180146
rect 193416 176730 193444 180118
rect 193404 176724 193456 176730
rect 193404 176666 193456 176672
rect 193876 161474 193904 180118
rect 194612 175642 194640 180118
rect 194888 176066 194916 180118
rect 195440 177410 195468 180118
rect 195428 177404 195480 177410
rect 195428 177346 195480 177352
rect 194704 176038 194916 176066
rect 194600 175636 194652 175642
rect 194600 175578 194652 175584
rect 193600 161446 193904 161474
rect 193312 4820 193364 4826
rect 193312 4762 193364 4768
rect 193220 4752 193272 4758
rect 193220 4694 193272 4700
rect 192024 3256 192076 3262
rect 192024 3198 192076 3204
rect 192036 480 192064 3198
rect 193232 480 193260 4694
rect 193600 3466 193628 161446
rect 194704 155242 194732 176038
rect 194784 175636 194836 175642
rect 194784 175578 194836 175584
rect 194692 155236 194744 155242
rect 194692 155178 194744 155184
rect 194416 7676 194468 7682
rect 194416 7618 194468 7624
rect 193588 3460 193640 3466
rect 193588 3402 193640 3408
rect 194428 480 194456 7618
rect 194796 4894 194824 175578
rect 195992 4962 196020 180118
rect 196452 161474 196480 180118
rect 197464 174570 197492 180118
rect 196084 161446 196480 161474
rect 197372 174542 197492 174570
rect 197556 180118 197846 180146
rect 198016 180118 198398 180146
rect 198752 180118 198858 180146
rect 198936 180118 199410 180146
rect 199580 180118 199962 180146
rect 200132 180118 200422 180146
rect 200592 180118 200974 180146
rect 201144 180118 201434 180146
rect 201604 180118 201986 180146
rect 202156 180118 202538 180146
rect 202892 180118 202998 180146
rect 203076 180118 203550 180146
rect 203720 180118 204010 180146
rect 204364 180118 204562 180146
rect 204824 180118 205114 180146
rect 205192 180118 205574 180146
rect 205652 180118 206126 180146
rect 206204 180118 206586 180146
rect 207032 180118 207138 180146
rect 207308 180118 207690 180146
rect 207768 180118 208150 180146
rect 208412 180118 208702 180146
rect 208780 180118 209162 180146
rect 209240 180118 209714 180146
rect 209792 180118 210266 180146
rect 210344 180118 210726 180146
rect 211278 180118 211384 180146
rect 196084 153882 196112 161446
rect 196072 153876 196124 153882
rect 196072 153818 196124 153824
rect 196808 7608 196860 7614
rect 196808 7550 196860 7556
rect 195980 4956 196032 4962
rect 195980 4898 196032 4904
rect 194784 4888 194836 4894
rect 194784 4830 194836 4836
rect 195612 3460 195664 3466
rect 195612 3402 195664 3408
rect 195624 480 195652 3402
rect 196820 480 196848 7550
rect 197372 3369 197400 174542
rect 197556 161474 197584 180118
rect 198016 171834 198044 180118
rect 198004 171828 198056 171834
rect 198004 171770 198056 171776
rect 197464 161446 197584 161474
rect 197464 5030 197492 161446
rect 197912 13116 197964 13122
rect 197912 13058 197964 13064
rect 197452 5024 197504 5030
rect 197452 4966 197504 4972
rect 197358 3360 197414 3369
rect 197358 3295 197414 3304
rect 197924 480 197952 13058
rect 198752 3534 198780 180118
rect 198936 170406 198964 180118
rect 198924 170400 198976 170406
rect 198924 170342 198976 170348
rect 199580 161474 199608 180118
rect 199028 161446 199608 161474
rect 199028 152522 199056 161446
rect 199016 152516 199068 152522
rect 199016 152458 199068 152464
rect 200132 3602 200160 180118
rect 200212 175636 200264 175642
rect 200212 175578 200264 175584
rect 200224 151094 200252 175578
rect 200592 169046 200620 180118
rect 201144 175642 201172 180118
rect 201500 177336 201552 177342
rect 201500 177278 201552 177284
rect 201132 175636 201184 175642
rect 201132 175578 201184 175584
rect 200580 169040 200632 169046
rect 200580 168982 200632 168988
rect 200212 151088 200264 151094
rect 200212 151030 200264 151036
rect 201512 11830 201540 177278
rect 201500 11824 201552 11830
rect 201500 11766 201552 11772
rect 200304 8968 200356 8974
rect 200304 8910 200356 8916
rect 200120 3596 200172 3602
rect 200120 3538 200172 3544
rect 198740 3528 198792 3534
rect 198740 3470 198792 3476
rect 199108 3528 199160 3534
rect 199108 3470 199160 3476
rect 199120 480 199148 3470
rect 200316 480 200344 8910
rect 201604 3670 201632 180118
rect 202156 167686 202184 180118
rect 202892 174554 202920 180118
rect 202880 174548 202932 174554
rect 202880 174490 202932 174496
rect 202144 167680 202196 167686
rect 202144 167622 202196 167628
rect 202696 11824 202748 11830
rect 202696 11766 202748 11772
rect 201684 10532 201736 10538
rect 201684 10474 201736 10480
rect 201592 3664 201644 3670
rect 201592 3606 201644 3612
rect 201696 3482 201724 10474
rect 201512 3454 201724 3482
rect 201512 480 201540 3454
rect 202708 480 202736 11766
rect 203076 3738 203104 180118
rect 203720 177682 203748 180118
rect 203708 177676 203760 177682
rect 203708 177618 203760 177624
rect 204260 171284 204312 171290
rect 204260 171226 204312 171232
rect 203892 6316 203944 6322
rect 203892 6258 203944 6264
rect 203064 3732 203116 3738
rect 203064 3674 203116 3680
rect 203904 480 203932 6258
rect 204272 3806 204300 171226
rect 204364 148374 204392 180118
rect 204824 171290 204852 180118
rect 204812 171284 204864 171290
rect 204812 171226 204864 171232
rect 205192 166326 205220 180118
rect 205652 173194 205680 180118
rect 206204 175658 206232 180118
rect 206284 177404 206336 177410
rect 206284 177346 206336 177352
rect 205744 175630 206232 175658
rect 205640 173188 205692 173194
rect 205640 173130 205692 173136
rect 205180 166320 205232 166326
rect 205180 166262 205232 166268
rect 204352 148368 204404 148374
rect 204352 148310 204404 148316
rect 205744 3874 205772 175630
rect 206296 161474 206324 177346
rect 207032 174622 207060 180118
rect 207204 175636 207256 175642
rect 207204 175578 207256 175584
rect 207020 174616 207072 174622
rect 207020 174558 207072 174564
rect 205836 161446 206324 161474
rect 205836 16574 205864 161446
rect 205836 16546 206232 16574
rect 205732 3868 205784 3874
rect 205732 3810 205784 3816
rect 204260 3800 204312 3806
rect 204260 3742 204312 3748
rect 205088 3120 205140 3126
rect 205088 3062 205140 3068
rect 205100 480 205128 3062
rect 206204 480 206232 16546
rect 207112 10328 207164 10334
rect 207112 10270 207164 10276
rect 190798 354 190910 480
rect 190472 326 190910 354
rect 190798 -960 190910 326
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207124 354 207152 10270
rect 207216 3942 207244 175578
rect 207308 164898 207336 180118
rect 207768 175642 207796 180118
rect 207756 175636 207808 175642
rect 207756 175578 207808 175584
rect 208412 173262 208440 180118
rect 208780 175658 208808 180118
rect 208504 175630 208808 175658
rect 208400 173256 208452 173262
rect 208400 173198 208452 173204
rect 207296 164892 207348 164898
rect 207296 164834 207348 164840
rect 208504 163538 208532 175630
rect 209240 171714 209268 180118
rect 209320 177676 209372 177682
rect 209320 177618 209372 177624
rect 208596 171686 209268 171714
rect 208492 163532 208544 163538
rect 208492 163474 208544 163480
rect 208596 4078 208624 171686
rect 209332 161474 209360 177618
rect 209792 171902 209820 180118
rect 210344 175658 210372 180118
rect 209884 175630 210372 175658
rect 209780 171896 209832 171902
rect 209780 171838 209832 171844
rect 209056 161446 209360 161474
rect 209056 10538 209084 161446
rect 209884 11762 209912 175630
rect 209964 172032 210016 172038
rect 209964 171974 210016 171980
rect 209976 16574 210004 171974
rect 209976 16546 211016 16574
rect 209872 11756 209924 11762
rect 209872 11698 209924 11704
rect 209044 10532 209096 10538
rect 209044 10474 209096 10480
rect 208584 4072 208636 4078
rect 208584 4014 208636 4020
rect 207204 3936 207256 3942
rect 207204 3878 207256 3884
rect 209780 3732 209832 3738
rect 209780 3674 209832 3680
rect 208584 3664 208636 3670
rect 208584 3606 208636 3612
rect 208596 480 208624 3606
rect 209792 480 209820 3674
rect 210988 480 211016 16546
rect 211356 4010 211384 180118
rect 211448 180118 211738 180146
rect 211908 180118 212290 180146
rect 212552 180118 212842 180146
rect 212920 180118 213302 180146
rect 213380 180118 213854 180146
rect 214024 180118 214314 180146
rect 214484 180118 214866 180146
rect 215312 180118 215418 180146
rect 215588 180118 215878 180146
rect 215956 180118 216430 180146
rect 216784 180118 216890 180146
rect 217152 180118 217442 180146
rect 217520 180118 217994 180146
rect 218164 180118 218454 180146
rect 218624 180118 219006 180146
rect 219466 180118 219572 180146
rect 211448 177614 211476 180118
rect 211436 177608 211488 177614
rect 211436 177550 211488 177556
rect 211908 162178 211936 180118
rect 211896 162172 211948 162178
rect 211896 162114 211948 162120
rect 212552 4146 212580 180118
rect 212920 175658 212948 180118
rect 212644 175630 212948 175658
rect 212644 5098 212672 175630
rect 213380 161474 213408 180118
rect 214024 177478 214052 180118
rect 214012 177472 214064 177478
rect 214012 177414 214064 177420
rect 214484 161474 214512 180118
rect 214564 177472 214616 177478
rect 214564 177414 214616 177420
rect 212736 161446 213408 161474
rect 214116 161446 214512 161474
rect 212736 160750 212764 161446
rect 212724 160744 212776 160750
rect 212724 160686 212776 160692
rect 214116 5166 214144 161446
rect 214576 6322 214604 177414
rect 215312 175930 215340 180118
rect 215312 175902 215432 175930
rect 215300 175636 215352 175642
rect 215300 175578 215352 175584
rect 214564 6316 214616 6322
rect 214564 6258 214616 6264
rect 214472 6248 214524 6254
rect 214472 6190 214524 6196
rect 214104 5160 214156 5166
rect 214104 5102 214156 5108
rect 212632 5092 212684 5098
rect 212632 5034 212684 5040
rect 212540 4140 212592 4146
rect 212540 4082 212592 4088
rect 211344 4004 211396 4010
rect 211344 3946 211396 3952
rect 213368 3868 213420 3874
rect 213368 3810 213420 3816
rect 212172 3800 212224 3806
rect 212172 3742 212224 3748
rect 212184 480 212212 3742
rect 213380 480 213408 3810
rect 214484 480 214512 6190
rect 215312 3398 215340 175578
rect 215404 171134 215432 175902
rect 215588 175642 215616 180118
rect 215576 175636 215628 175642
rect 215576 175578 215628 175584
rect 215404 171106 215524 171134
rect 215496 159390 215524 171106
rect 215956 161474 215984 180118
rect 215588 161446 215984 161474
rect 215484 159384 215536 159390
rect 215484 159326 215536 159332
rect 215588 5234 215616 161446
rect 216784 158030 216812 180118
rect 217152 177546 217180 180118
rect 217140 177540 217192 177546
rect 217140 177482 217192 177488
rect 217520 175658 217548 180118
rect 217600 176928 217652 176934
rect 217600 176870 217652 176876
rect 216968 175630 217548 175658
rect 216772 158024 216824 158030
rect 216772 157966 216824 157972
rect 216968 6186 216996 175630
rect 217612 161474 217640 176870
rect 218060 175636 218112 175642
rect 218060 175578 218112 175584
rect 217336 161446 217640 161474
rect 217336 7682 217364 161446
rect 218072 16574 218100 175578
rect 218164 170474 218192 180118
rect 218624 175642 218652 180118
rect 218612 175636 218664 175642
rect 218612 175578 218664 175584
rect 218152 170468 218204 170474
rect 218152 170410 218204 170416
rect 218072 16546 218192 16574
rect 217324 7676 217376 7682
rect 217324 7618 217376 7624
rect 216956 6180 217008 6186
rect 216956 6122 217008 6128
rect 215576 5228 215628 5234
rect 215576 5170 215628 5176
rect 218060 4888 218112 4894
rect 218060 4830 218112 4836
rect 215668 4004 215720 4010
rect 215668 3946 215720 3952
rect 215300 3392 215352 3398
rect 215300 3334 215352 3340
rect 215680 480 215708 3946
rect 216864 3936 216916 3942
rect 216864 3878 216916 3884
rect 216876 480 216904 3878
rect 218072 480 218100 4830
rect 218164 3330 218192 16546
rect 219544 5302 219572 180118
rect 219636 180118 220018 180146
rect 220188 180118 220570 180146
rect 220924 180118 221030 180146
rect 221200 180118 221582 180146
rect 221660 180118 222042 180146
rect 222212 180118 222594 180146
rect 222764 180118 223146 180146
rect 223606 180118 223712 180146
rect 219636 169114 219664 180118
rect 219624 169108 219676 169114
rect 219624 169050 219676 169056
rect 220188 161474 220216 180118
rect 219728 161446 220216 161474
rect 219532 5296 219584 5302
rect 219532 5238 219584 5244
rect 219256 4140 219308 4146
rect 219256 4082 219308 4088
rect 218152 3324 218204 3330
rect 218152 3266 218204 3272
rect 219268 480 219296 4082
rect 219728 3262 219756 161446
rect 220924 4826 220952 180118
rect 221200 176934 221228 180118
rect 221188 176928 221240 176934
rect 221188 176870 221240 176876
rect 221660 161474 221688 180118
rect 221108 161446 221688 161474
rect 220912 4820 220964 4826
rect 220912 4762 220964 4768
rect 220452 4072 220504 4078
rect 220452 4014 220504 4020
rect 219716 3256 219768 3262
rect 219716 3198 219768 3204
rect 220464 480 220492 4014
rect 221108 3466 221136 161446
rect 222212 7614 222240 180118
rect 222764 161474 222792 180118
rect 223684 175624 223712 180118
rect 223776 180118 224158 180146
rect 224236 180118 224618 180146
rect 224972 180118 225170 180146
rect 225432 180118 225722 180146
rect 225800 180118 226182 180146
rect 226536 180118 226734 180146
rect 226904 180118 227286 180146
rect 227746 180118 227852 180146
rect 223776 175982 223804 180118
rect 223764 175976 223816 175982
rect 223764 175918 223816 175924
rect 222304 161446 222792 161474
rect 223592 175596 223712 175624
rect 222304 13122 222332 161446
rect 222292 13116 222344 13122
rect 222292 13058 222344 13064
rect 222200 7608 222252 7614
rect 222200 7550 222252 7556
rect 223592 3534 223620 175596
rect 224236 161474 224264 180118
rect 224972 177682 225000 180118
rect 224960 177676 225012 177682
rect 224960 177618 225012 177624
rect 225432 177342 225460 180118
rect 225800 177478 225828 180118
rect 225788 177472 225840 177478
rect 225788 177414 225840 177420
rect 225420 177336 225472 177342
rect 225420 177278 225472 177284
rect 226340 176996 226392 177002
rect 226340 176938 226392 176944
rect 226352 172038 226380 176938
rect 226340 172032 226392 172038
rect 226340 171974 226392 171980
rect 223684 161446 224264 161474
rect 223684 8974 223712 161446
rect 223672 8968 223724 8974
rect 223672 8910 223724 8916
rect 223580 3528 223632 3534
rect 223580 3470 223632 3476
rect 223948 3528 224000 3534
rect 223948 3470 224000 3476
rect 221096 3460 221148 3466
rect 221096 3402 221148 3408
rect 222752 3392 222804 3398
rect 222752 3334 222804 3340
rect 221556 3188 221608 3194
rect 221556 3130 221608 3136
rect 221568 480 221596 3130
rect 222764 480 222792 3334
rect 223960 480 223988 3470
rect 225144 3324 225196 3330
rect 225144 3266 225196 3272
rect 225156 480 225184 3266
rect 226340 3256 226392 3262
rect 226340 3198 226392 3204
rect 226352 480 226380 3198
rect 226536 3126 226564 180118
rect 226904 177410 226932 180118
rect 226892 177404 226944 177410
rect 226892 177346 226944 177352
rect 227824 176730 227852 180118
rect 228008 180118 228298 180146
rect 228376 180118 228758 180146
rect 229204 180118 229310 180146
rect 229388 180118 229862 180146
rect 230032 180118 230322 180146
rect 230584 180118 230874 180146
rect 230952 180118 231334 180146
rect 231886 180118 231992 180146
rect 227904 177608 227956 177614
rect 227904 177550 227956 177556
rect 226984 176724 227036 176730
rect 226984 176666 227036 176672
rect 227812 176724 227864 176730
rect 227812 176666 227864 176672
rect 226996 10334 227024 176666
rect 227916 174298 227944 177550
rect 227732 174270 227944 174298
rect 226984 10328 227036 10334
rect 226984 10270 227036 10276
rect 227536 3732 227588 3738
rect 227536 3674 227588 3680
rect 226524 3120 226576 3126
rect 226524 3062 226576 3068
rect 227548 480 227576 3674
rect 227732 490 227760 174270
rect 228008 174162 228036 180118
rect 227824 174134 228036 174162
rect 227824 3602 227852 174134
rect 228376 161474 228404 180118
rect 229204 177002 229232 180118
rect 229192 176996 229244 177002
rect 229192 176938 229244 176944
rect 229192 175636 229244 175642
rect 229192 175578 229244 175584
rect 227916 161446 228404 161474
rect 227916 3670 227944 161446
rect 229204 3874 229232 175578
rect 229192 3868 229244 3874
rect 229192 3810 229244 3816
rect 229388 3806 229416 180118
rect 230032 175642 230060 180118
rect 230020 175636 230072 175642
rect 230020 175578 230072 175584
rect 230480 175636 230532 175642
rect 230480 175578 230532 175584
rect 230492 4010 230520 175578
rect 230584 6254 230612 180118
rect 230952 175642 230980 180118
rect 230940 175636 230992 175642
rect 230940 175578 230992 175584
rect 230572 6248 230624 6254
rect 230572 6190 230624 6196
rect 230480 4004 230532 4010
rect 230480 3946 230532 3952
rect 231964 3942 231992 180118
rect 232056 180118 232438 180146
rect 232608 180118 232898 180146
rect 233252 180118 233450 180146
rect 233620 180118 233910 180146
rect 234080 180118 234462 180146
rect 234632 180118 235014 180146
rect 235184 180118 235474 180146
rect 236026 180118 236132 180146
rect 232056 4894 232084 180118
rect 232608 161474 232636 180118
rect 232148 161446 232636 161474
rect 232044 4888 232096 4894
rect 232044 4830 232096 4836
rect 232148 4146 232176 161446
rect 232136 4140 232188 4146
rect 232136 4082 232188 4088
rect 233252 4078 233280 180118
rect 233332 175636 233384 175642
rect 233332 175578 233384 175584
rect 233240 4072 233292 4078
rect 233240 4014 233292 4020
rect 231952 3936 232004 3942
rect 231952 3878 232004 3884
rect 229376 3800 229428 3806
rect 229376 3742 229428 3748
rect 227904 3664 227956 3670
rect 227904 3606 227956 3612
rect 229836 3664 229888 3670
rect 229836 3606 229888 3612
rect 227812 3596 227864 3602
rect 227812 3538 227864 3544
rect 207358 354 207470 480
rect 207124 326 207470 354
rect 207358 -960 207470 326
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 227732 462 228312 490
rect 229848 480 229876 3606
rect 232228 3596 232280 3602
rect 232228 3538 232280 3544
rect 231032 3460 231084 3466
rect 231032 3402 231084 3408
rect 231044 480 231072 3402
rect 232240 480 232268 3538
rect 233344 3398 233372 175578
rect 233332 3392 233384 3398
rect 233332 3334 233384 3340
rect 233620 3194 233648 180118
rect 234080 175642 234108 180118
rect 234068 175636 234120 175642
rect 234068 175578 234120 175584
rect 234632 3534 234660 180118
rect 234712 176928 234764 176934
rect 234712 176870 234764 176876
rect 234620 3528 234672 3534
rect 234620 3470 234672 3476
rect 234724 3210 234752 176870
rect 235184 161474 235212 180118
rect 235264 176724 235316 176730
rect 235264 176666 235316 176672
rect 234816 161446 235212 161474
rect 234816 3330 234844 161446
rect 235276 3602 235304 176666
rect 236104 174706 236132 180118
rect 236012 174678 236132 174706
rect 236196 180118 236486 180146
rect 236656 180118 237038 180146
rect 237484 180118 237590 180146
rect 237668 180118 238050 180146
rect 238312 180118 238602 180146
rect 238864 180118 239062 180146
rect 239140 180118 239614 180146
rect 240166 180118 240272 180146
rect 235264 3596 235316 3602
rect 235264 3538 235316 3544
rect 234804 3324 234856 3330
rect 234804 3266 234856 3272
rect 236012 3262 236040 174678
rect 236092 174004 236144 174010
rect 236092 173946 236144 173952
rect 236000 3256 236052 3262
rect 233608 3188 233660 3194
rect 234724 3182 235856 3210
rect 236000 3198 236052 3204
rect 236104 3210 236132 173946
rect 236196 3738 236224 180118
rect 236656 177614 236684 180118
rect 236644 177608 236696 177614
rect 236644 177550 236696 177556
rect 236276 176860 236328 176866
rect 236276 176802 236328 176808
rect 236288 174010 236316 176802
rect 236276 174004 236328 174010
rect 236276 173946 236328 173952
rect 236184 3732 236236 3738
rect 236184 3674 236236 3680
rect 237484 3670 237512 180118
rect 237472 3664 237524 3670
rect 237472 3606 237524 3612
rect 237668 3466 237696 180118
rect 238024 176996 238076 177002
rect 238024 176938 238076 176944
rect 237656 3460 237708 3466
rect 237656 3402 237708 3408
rect 236104 3182 236592 3210
rect 233608 3130 233660 3136
rect 234620 3052 234672 3058
rect 234620 2994 234672 3000
rect 233424 2916 233476 2922
rect 233424 2858 233476 2864
rect 233436 480 233464 2858
rect 234632 480 234660 2994
rect 235828 480 235856 3182
rect 228284 354 228312 462
rect 228702 354 228814 480
rect 228284 326 228814 354
rect 228702 -960 228814 326
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236564 354 236592 3182
rect 238036 2922 238064 176938
rect 238312 176730 238340 180118
rect 238864 177002 238892 180118
rect 238852 176996 238904 177002
rect 238852 176938 238904 176944
rect 238300 176724 238352 176730
rect 238300 176666 238352 176672
rect 239140 161474 239168 180118
rect 240244 176934 240272 180118
rect 240336 180118 240626 180146
rect 240704 180118 241178 180146
rect 241532 180118 241638 180146
rect 241808 180118 242190 180146
rect 242360 180118 242742 180146
rect 243004 180118 243202 180146
rect 243464 180118 243754 180146
rect 244108 180118 244214 180146
rect 244766 180118 244872 180146
rect 240232 176928 240284 176934
rect 240232 176870 240284 176876
rect 240336 176866 240364 180118
rect 240324 176860 240376 176866
rect 240324 176802 240376 176808
rect 240704 161474 240732 180118
rect 241532 176730 241560 180118
rect 240784 176724 240836 176730
rect 240784 176666 240836 176672
rect 241520 176724 241572 176730
rect 241520 176666 241572 176672
rect 238956 161446 239168 161474
rect 240336 161446 240732 161474
rect 238116 3732 238168 3738
rect 238116 3674 238168 3680
rect 238024 2916 238076 2922
rect 238024 2858 238076 2864
rect 238128 480 238156 3674
rect 238956 3058 238984 161446
rect 240336 3738 240364 161446
rect 240324 3732 240376 3738
rect 240324 3674 240376 3680
rect 240796 3534 240824 176666
rect 241704 175636 241756 175642
rect 241704 175578 241756 175584
rect 239312 3528 239364 3534
rect 239312 3470 239364 3476
rect 240784 3528 240836 3534
rect 240784 3470 240836 3476
rect 238944 3052 238996 3058
rect 238944 2994 238996 3000
rect 239324 480 239352 3470
rect 240508 3460 240560 3466
rect 240508 3402 240560 3408
rect 240520 480 240548 3402
rect 241716 480 241744 175578
rect 241808 3466 241836 180118
rect 242360 175642 242388 180118
rect 242348 175636 242400 175642
rect 242348 175578 242400 175584
rect 242900 175636 242952 175642
rect 242900 175578 242952 175584
rect 242912 11762 242940 175578
rect 242900 11756 242952 11762
rect 242900 11698 242952 11704
rect 243004 6914 243032 180118
rect 243464 175642 243492 180118
rect 244108 176746 244136 180118
rect 244108 176718 244320 176746
rect 244844 176730 244872 180118
rect 244936 180118 245318 180146
rect 245778 180118 246160 180146
rect 243452 175636 243504 175642
rect 243452 175578 243504 175584
rect 244096 11756 244148 11762
rect 244096 11698 244148 11704
rect 242912 6886 243032 6914
rect 241796 3460 241848 3466
rect 241796 3402 241848 3408
rect 242912 480 242940 6886
rect 244108 480 244136 11698
rect 244292 3482 244320 176718
rect 244832 176724 244884 176730
rect 244832 176666 244884 176672
rect 244936 161474 244964 180118
rect 246132 177274 246160 180118
rect 246224 180118 246330 180146
rect 246408 180118 246790 180146
rect 247342 180118 247632 180146
rect 247894 180118 248184 180146
rect 246224 177410 246252 180118
rect 246212 177404 246264 177410
rect 246212 177346 246264 177352
rect 246120 177268 246172 177274
rect 246120 177210 246172 177216
rect 246408 176882 246436 180118
rect 247604 177342 247632 180118
rect 248156 177478 248184 180118
rect 248248 180118 248354 180146
rect 248616 180118 248906 180146
rect 248984 180118 249366 180146
rect 249812 180118 249918 180146
rect 249996 180118 250470 180146
rect 250548 180118 250930 180146
rect 251192 180118 251482 180146
rect 251942 180118 252232 180146
rect 248248 177546 248276 180118
rect 248236 177540 248288 177546
rect 248236 177482 248288 177488
rect 248144 177472 248196 177478
rect 248144 177414 248196 177420
rect 247592 177336 247644 177342
rect 247592 177278 247644 177284
rect 248420 177268 248472 177274
rect 248420 177210 248472 177216
rect 244384 161446 244964 161474
rect 245672 176854 246436 176882
rect 244384 3602 244412 161446
rect 245672 3670 245700 176854
rect 245752 176724 245804 176730
rect 245752 176666 245804 176672
rect 245764 16574 245792 176666
rect 245764 16546 245976 16574
rect 245660 3664 245712 3670
rect 245660 3606 245712 3612
rect 244372 3596 244424 3602
rect 244372 3538 244424 3544
rect 244292 3454 245240 3482
rect 245212 480 245240 3454
rect 236982 354 237094 480
rect 236564 326 237094 354
rect 236982 -960 237094 326
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 245948 354 245976 16546
rect 247592 3596 247644 3602
rect 247592 3538 247644 3544
rect 247604 480 247632 3538
rect 246366 354 246478 480
rect 245948 326 246478 354
rect 246366 -960 246478 326
rect 247562 -960 247674 480
rect 248432 354 248460 177210
rect 248512 171828 248564 171834
rect 248512 171770 248564 171776
rect 248524 3330 248552 171770
rect 248512 3324 248564 3330
rect 248512 3266 248564 3272
rect 248616 3058 248644 180118
rect 248984 171834 249012 180118
rect 249812 175658 249840 180118
rect 249812 175630 249932 175658
rect 249800 175568 249852 175574
rect 249800 175510 249852 175516
rect 248972 171828 249024 171834
rect 248972 171770 249024 171776
rect 249812 3482 249840 175510
rect 249904 3602 249932 175630
rect 249996 5114 250024 180118
rect 250076 177404 250128 177410
rect 250076 177346 250128 177352
rect 250088 175574 250116 177346
rect 250076 175568 250128 175574
rect 250076 175510 250128 175516
rect 250548 161474 250576 180118
rect 250088 161446 250576 161474
rect 250088 6254 250116 161446
rect 250076 6248 250128 6254
rect 250076 6190 250128 6196
rect 249996 5086 250116 5114
rect 249892 3596 249944 3602
rect 249892 3538 249944 3544
rect 249812 3454 250024 3482
rect 250088 3466 250116 5086
rect 251192 4146 251220 180118
rect 251824 177540 251876 177546
rect 251824 177482 251876 177488
rect 251272 177336 251324 177342
rect 251272 177278 251324 177284
rect 251284 16574 251312 177278
rect 251284 16546 251772 16574
rect 251180 4140 251232 4146
rect 251180 4082 251232 4088
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 248604 3052 248656 3058
rect 248604 2994 248656 3000
rect 249996 480 250024 3454
rect 250076 3460 250128 3466
rect 250076 3402 250128 3408
rect 251192 480 251220 3606
rect 251744 3482 251772 16546
rect 251836 3602 251864 177482
rect 252204 177410 252232 180118
rect 252388 180118 252494 180146
rect 252664 180118 253046 180146
rect 253124 180118 253506 180146
rect 254058 180118 254164 180146
rect 252192 177404 252244 177410
rect 252192 177346 252244 177352
rect 252388 177342 252416 180118
rect 252560 177472 252612 177478
rect 252560 177414 252612 177420
rect 252376 177336 252428 177342
rect 252376 177278 252428 177284
rect 251824 3596 251876 3602
rect 251824 3538 251876 3544
rect 252572 3482 252600 177414
rect 252664 3942 252692 180118
rect 253124 161474 253152 180118
rect 254136 175658 254164 180118
rect 253940 175636 253992 175642
rect 253940 175578 253992 175584
rect 254044 175630 254164 175658
rect 254228 180118 254518 180146
rect 254688 180118 255070 180146
rect 255424 180118 255622 180146
rect 255700 180118 256082 180146
rect 256344 180118 256634 180146
rect 256712 180118 257094 180146
rect 257264 180118 257646 180146
rect 258092 180118 258198 180146
rect 258368 180118 258658 180146
rect 258920 180118 259210 180146
rect 259472 180118 259762 180146
rect 259840 180118 260222 180146
rect 260392 180118 260774 180146
rect 260852 180118 261234 180146
rect 261786 180118 262168 180146
rect 252756 161446 253152 161474
rect 252652 3936 252704 3942
rect 252652 3878 252704 3884
rect 252756 3874 252784 161446
rect 252744 3868 252796 3874
rect 252744 3810 252796 3816
rect 253952 3806 253980 175578
rect 254044 13122 254072 175630
rect 254228 161474 254256 180118
rect 254688 175642 254716 180118
rect 254676 175636 254728 175642
rect 254676 175578 254728 175584
rect 255320 175636 255372 175642
rect 255320 175578 255372 175584
rect 254136 161446 254256 161474
rect 254136 29646 254164 161446
rect 254124 29640 254176 29646
rect 254124 29582 254176 29588
rect 254032 13116 254084 13122
rect 254032 13058 254084 13064
rect 253940 3800 253992 3806
rect 253940 3742 253992 3748
rect 255332 3738 255360 175578
rect 255424 4894 255452 180118
rect 255700 161474 255728 180118
rect 256344 175642 256372 180118
rect 256332 175636 256384 175642
rect 256332 175578 256384 175584
rect 255516 161446 255728 161474
rect 255516 6186 255544 161446
rect 256712 7682 256740 180118
rect 257264 161474 257292 180118
rect 256804 161446 257292 161474
rect 256804 18834 256832 161446
rect 256792 18828 256844 18834
rect 256792 18770 256844 18776
rect 256700 7676 256752 7682
rect 256700 7618 256752 7624
rect 255504 6180 255556 6186
rect 255504 6122 255556 6128
rect 255412 4888 255464 4894
rect 255412 4830 255464 4836
rect 255320 3732 255372 3738
rect 255320 3674 255372 3680
rect 258092 3670 258120 180118
rect 258264 174140 258316 174146
rect 258264 174082 258316 174088
rect 258276 4826 258304 174082
rect 258368 9042 258396 180118
rect 258920 174146 258948 180118
rect 258908 174140 258960 174146
rect 258908 174082 258960 174088
rect 258356 9036 258408 9042
rect 258356 8978 258408 8984
rect 258264 4820 258316 4826
rect 258264 4762 258316 4768
rect 258080 3664 258132 3670
rect 258080 3606 258132 3612
rect 259472 3602 259500 180118
rect 259552 175636 259604 175642
rect 259552 175578 259604 175584
rect 259564 7614 259592 175578
rect 259840 161474 259868 180118
rect 260392 175642 260420 180118
rect 260380 175636 260432 175642
rect 260380 175578 260432 175584
rect 259656 161446 259868 161474
rect 259656 11898 259684 161446
rect 259644 11892 259696 11898
rect 259644 11834 259696 11840
rect 259552 7608 259604 7614
rect 259552 7550 259604 7556
rect 260656 6248 260708 6254
rect 260656 6190 260708 6196
rect 254676 3596 254728 3602
rect 254676 3538 254728 3544
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 251744 3454 252416 3482
rect 252572 3454 253520 3482
rect 252388 480 252416 3454
rect 253492 480 253520 3454
rect 254688 480 254716 3538
rect 258264 3528 258316 3534
rect 258264 3470 258316 3476
rect 257068 3324 257120 3330
rect 257068 3266 257120 3272
rect 255872 3052 255924 3058
rect 255872 2994 255924 3000
rect 255884 480 255912 2994
rect 257080 480 257108 3266
rect 258276 480 258304 3470
rect 259460 3460 259512 3466
rect 259460 3402 259512 3408
rect 259472 480 259500 3402
rect 260668 480 260696 6190
rect 260852 3534 260880 180118
rect 262140 176934 262168 180118
rect 262232 180118 262338 180146
rect 262416 180118 262798 180146
rect 262876 180118 263350 180146
rect 263810 180118 263916 180146
rect 264362 180118 264560 180146
rect 262232 177546 262260 180118
rect 262220 177540 262272 177546
rect 262220 177482 262272 177488
rect 262220 177404 262272 177410
rect 262220 177346 262272 177352
rect 262128 176928 262180 176934
rect 262128 176870 262180 176876
rect 262232 16574 262260 177346
rect 262232 16546 262352 16574
rect 261760 4140 261812 4146
rect 261760 4082 261812 4088
rect 260840 3528 260892 3534
rect 260840 3470 260892 3476
rect 261772 480 261800 4082
rect 262324 490 262352 16546
rect 262416 3466 262444 180118
rect 262876 161474 262904 180118
rect 263600 177336 263652 177342
rect 263600 177278 263652 177284
rect 262508 161446 262904 161474
rect 262508 10470 262536 161446
rect 262496 10464 262548 10470
rect 262496 10406 262548 10412
rect 263612 6914 263640 177278
rect 263692 175636 263744 175642
rect 263692 175578 263744 175584
rect 263704 8974 263732 175578
rect 263888 161474 263916 180118
rect 264532 177410 264560 180118
rect 264624 180118 264914 180146
rect 265268 180118 265374 180146
rect 265452 180118 265926 180146
rect 266386 180118 266492 180146
rect 264520 177404 264572 177410
rect 264520 177346 264572 177352
rect 264624 175642 264652 180118
rect 265268 177546 265296 180118
rect 265256 177540 265308 177546
rect 265256 177482 265308 177488
rect 264612 175636 264664 175642
rect 264612 175578 264664 175584
rect 265452 161474 265480 180118
rect 266464 174434 266492 180118
rect 263796 161446 263916 161474
rect 264992 161446 265480 161474
rect 266372 174406 266492 174434
rect 266556 180118 266938 180146
rect 267016 180118 267490 180146
rect 267752 180118 267950 180146
rect 268028 180118 268502 180146
rect 268672 180118 268962 180146
rect 269224 180118 269514 180146
rect 269776 180118 270066 180146
rect 270526 180118 270632 180146
rect 263796 10402 263824 161446
rect 264992 24138 265020 161446
rect 264980 24132 265032 24138
rect 264980 24074 265032 24080
rect 266372 17270 266400 174406
rect 266556 174298 266584 180118
rect 266464 174270 266584 174298
rect 266360 17264 266412 17270
rect 266360 17206 266412 17212
rect 266464 13190 266492 174270
rect 267016 161474 267044 180118
rect 266556 161446 267044 161474
rect 266556 25566 266584 161446
rect 266544 25560 266596 25566
rect 266544 25502 266596 25508
rect 267752 22778 267780 180118
rect 267832 175636 267884 175642
rect 267832 175578 267884 175584
rect 267844 26926 267872 175578
rect 268028 29646 268056 180118
rect 268672 175642 268700 180118
rect 268660 175636 268712 175642
rect 268660 175578 268712 175584
rect 269120 175636 269172 175642
rect 269120 175578 269172 175584
rect 267924 29640 267976 29646
rect 267924 29582 267976 29588
rect 268016 29640 268068 29646
rect 268016 29582 268068 29588
rect 267832 26920 267884 26926
rect 267832 26862 267884 26868
rect 267740 22772 267792 22778
rect 267740 22714 267792 22720
rect 267936 16574 267964 29582
rect 267936 16546 268424 16574
rect 266452 13184 266504 13190
rect 266452 13126 266504 13132
rect 267740 13116 267792 13122
rect 267740 13058 267792 13064
rect 263784 10396 263836 10402
rect 263784 10338 263836 10344
rect 263692 8968 263744 8974
rect 263692 8910 263744 8916
rect 263612 6886 264192 6914
rect 262404 3460 262456 3466
rect 262404 3402 262456 3408
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262324 462 262536 490
rect 264164 480 264192 6886
rect 265348 3936 265400 3942
rect 265348 3878 265400 3884
rect 265360 480 265388 3878
rect 266544 3868 266596 3874
rect 266544 3810 266596 3816
rect 266556 480 266584 3810
rect 267752 480 267780 13058
rect 262508 354 262536 462
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 269132 6254 269160 175578
rect 269224 13122 269252 180118
rect 269672 176928 269724 176934
rect 269672 176870 269724 176876
rect 269684 171134 269712 176870
rect 269776 175642 269804 180118
rect 270604 175658 270632 180118
rect 269764 175636 269816 175642
rect 269764 175578 269816 175584
rect 270512 175630 270632 175658
rect 270696 180118 271078 180146
rect 271156 180118 271538 180146
rect 271892 180118 272090 180146
rect 272642 180118 273024 180146
rect 273102 180118 273208 180146
rect 269684 171106 269804 171134
rect 269212 13116 269264 13122
rect 269212 13058 269264 13064
rect 269120 6248 269172 6254
rect 269120 6190 269172 6196
rect 269776 4962 269804 171106
rect 270512 31074 270540 175630
rect 270696 175522 270724 180118
rect 270604 175494 270724 175522
rect 270500 31068 270552 31074
rect 270500 31010 270552 31016
rect 270604 14550 270632 175494
rect 271156 161474 271184 180118
rect 270696 161446 271184 161474
rect 270696 21486 270724 161446
rect 271892 35222 271920 180118
rect 272996 176730 273024 180118
rect 273180 176934 273208 180118
rect 273364 180118 273654 180146
rect 273824 180118 274114 180146
rect 274666 180118 274772 180146
rect 273168 176928 273220 176934
rect 273168 176870 273220 176876
rect 272984 176724 273036 176730
rect 272984 176666 273036 176672
rect 273260 171828 273312 171834
rect 273260 171770 273312 171776
rect 271880 35216 271932 35222
rect 271880 35158 271932 35164
rect 270684 21480 270736 21486
rect 270684 21422 270736 21428
rect 270592 14544 270644 14550
rect 270592 14486 270644 14492
rect 273272 11830 273300 171770
rect 273364 37942 273392 180118
rect 273824 171834 273852 180118
rect 273904 176724 273956 176730
rect 273904 176666 273956 176672
rect 273812 171828 273864 171834
rect 273812 171770 273864 171776
rect 273352 37936 273404 37942
rect 273352 37878 273404 37884
rect 273916 15978 273944 176666
rect 274744 166994 274772 180118
rect 274652 166966 274772 166994
rect 274928 180118 275218 180146
rect 275678 180118 275968 180146
rect 273904 15972 273956 15978
rect 273904 15914 273956 15920
rect 273260 11824 273312 11830
rect 273260 11766 273312 11772
rect 274652 10334 274680 166966
rect 274928 161474 274956 180118
rect 275940 175982 275968 180118
rect 276032 180118 276230 180146
rect 276308 180118 276690 180146
rect 276952 180118 277242 180146
rect 277412 180118 277794 180146
rect 277872 180118 278254 180146
rect 278806 180118 279096 180146
rect 275928 175976 275980 175982
rect 275928 175918 275980 175924
rect 274744 161446 274956 161474
rect 274744 14482 274772 161446
rect 276032 16574 276060 180118
rect 276112 167068 276164 167074
rect 276112 167010 276164 167016
rect 276124 18698 276152 167010
rect 276308 39370 276336 180118
rect 276952 167074 276980 180118
rect 276940 167068 276992 167074
rect 276940 167010 276992 167016
rect 276296 39364 276348 39370
rect 276296 39306 276348 39312
rect 276204 18828 276256 18834
rect 276204 18770 276256 18776
rect 276112 18692 276164 18698
rect 276112 18634 276164 18640
rect 276032 16546 276152 16574
rect 274732 14476 274784 14482
rect 274732 14418 274784 14424
rect 274640 10328 274692 10334
rect 274640 10270 274692 10276
rect 274824 7676 274876 7682
rect 274824 7618 274876 7624
rect 272432 6180 272484 6186
rect 272432 6122 272484 6128
rect 269764 4956 269816 4962
rect 269764 4898 269816 4904
rect 271236 4888 271288 4894
rect 271236 4830 271288 4836
rect 270040 3800 270092 3806
rect 270040 3742 270092 3748
rect 270052 480 270080 3742
rect 271248 480 271276 4830
rect 272444 480 272472 6122
rect 273628 3732 273680 3738
rect 273628 3674 273680 3680
rect 273640 480 273668 3674
rect 274836 480 274864 7618
rect 276124 6594 276152 16546
rect 276112 6588 276164 6594
rect 276112 6530 276164 6536
rect 276216 3482 276244 18770
rect 277412 6526 277440 180118
rect 277872 161474 277900 180118
rect 278044 176928 278096 176934
rect 278044 176870 278096 176876
rect 277504 161446 277900 161474
rect 277504 40730 277532 161446
rect 277492 40724 277544 40730
rect 277492 40666 277544 40672
rect 278056 32502 278084 176870
rect 279068 176730 279096 180118
rect 279160 180118 279266 180146
rect 279344 180118 279818 180146
rect 280264 180118 280370 180146
rect 280448 180118 280830 180146
rect 280908 180118 281382 180146
rect 281736 180118 281842 180146
rect 281920 180118 282394 180146
rect 282946 180118 283052 180146
rect 283406 180118 283696 180146
rect 283958 180118 284248 180146
rect 279056 176724 279108 176730
rect 279056 176666 279108 176672
rect 279160 173194 279188 180118
rect 279148 173188 279200 173194
rect 279148 173130 279200 173136
rect 279344 161474 279372 180118
rect 280264 176654 280292 180118
rect 280264 176626 280384 176654
rect 280160 171828 280212 171834
rect 280160 171770 280212 171776
rect 278884 161446 279372 161474
rect 278884 46238 278912 161446
rect 278872 46232 278924 46238
rect 278872 46174 278924 46180
rect 278044 32496 278096 32502
rect 278044 32438 278096 32444
rect 278320 9036 278372 9042
rect 278320 8978 278372 8984
rect 277400 6520 277452 6526
rect 277400 6462 277452 6468
rect 277124 3664 277176 3670
rect 277124 3606 277176 3612
rect 276032 3454 276244 3482
rect 276032 480 276060 3454
rect 277136 480 277164 3606
rect 278332 480 278360 8978
rect 280172 6186 280200 171770
rect 280356 161474 280384 176626
rect 280448 171834 280476 180118
rect 280436 171828 280488 171834
rect 280436 171770 280488 171776
rect 280908 161474 280936 180118
rect 281736 177342 281764 180118
rect 281724 177336 281776 177342
rect 281724 177278 281776 177284
rect 281920 161474 281948 180118
rect 282184 177540 282236 177546
rect 282184 177482 282236 177488
rect 280264 161446 280384 161474
rect 280448 161446 280936 161474
rect 281552 161446 281948 161474
rect 280264 20058 280292 161446
rect 280448 123486 280476 161446
rect 280436 123480 280488 123486
rect 280436 123422 280488 123428
rect 280252 20052 280304 20058
rect 280252 19994 280304 20000
rect 281552 11762 281580 161446
rect 281632 11892 281684 11898
rect 281632 11834 281684 11840
rect 281540 11756 281592 11762
rect 281540 11698 281592 11704
rect 280160 6180 280212 6186
rect 280160 6122 280212 6128
rect 279516 4820 279568 4826
rect 279516 4762 279568 4768
rect 279528 480 279556 4762
rect 280712 3596 280764 3602
rect 280712 3538 280764 3544
rect 280724 480 280752 3538
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281644 354 281672 11834
rect 282196 9042 282224 177482
rect 282276 176724 282328 176730
rect 282276 176666 282328 176672
rect 282288 28286 282316 176666
rect 283024 161474 283052 180118
rect 283668 174554 283696 180118
rect 284220 177002 284248 180118
rect 284312 180118 284418 180146
rect 284680 180118 284970 180146
rect 285048 180118 285522 180146
rect 285982 180118 286272 180146
rect 284208 176996 284260 177002
rect 284208 176938 284260 176944
rect 284312 175624 284340 180118
rect 284312 175596 284432 175624
rect 284300 175500 284352 175506
rect 284300 175442 284352 175448
rect 283656 174548 283708 174554
rect 283656 174490 283708 174496
rect 282932 161446 283052 161474
rect 282276 28280 282328 28286
rect 282276 28222 282328 28228
rect 282932 15910 282960 161446
rect 282920 15904 282972 15910
rect 282920 15846 282972 15852
rect 282184 9036 282236 9042
rect 282184 8978 282236 8984
rect 283104 7608 283156 7614
rect 283104 7550 283156 7556
rect 283116 480 283144 7550
rect 284312 5234 284340 175442
rect 284404 21418 284432 175596
rect 284680 175506 284708 180118
rect 284668 175500 284720 175506
rect 284668 175442 284720 175448
rect 285048 161474 285076 180118
rect 286244 177478 286272 180118
rect 286336 180118 286534 180146
rect 286704 180118 286994 180146
rect 287164 180118 287546 180146
rect 287808 180118 288098 180146
rect 288452 180118 288558 180146
rect 288636 180118 289110 180146
rect 289280 180118 289570 180146
rect 290122 180118 290228 180146
rect 285680 177472 285732 177478
rect 285680 177414 285732 177420
rect 286232 177472 286284 177478
rect 286232 177414 286284 177420
rect 284496 161446 285076 161474
rect 284392 21412 284444 21418
rect 284392 21354 284444 21360
rect 284496 7682 284524 161446
rect 284484 7676 284536 7682
rect 284484 7618 284536 7624
rect 284300 5228 284352 5234
rect 284300 5170 284352 5176
rect 285404 4956 285456 4962
rect 285404 4898 285456 4904
rect 284300 3528 284352 3534
rect 284300 3470 284352 3476
rect 284312 480 284340 3470
rect 285416 480 285444 4898
rect 285692 3482 285720 177414
rect 286336 175624 286364 180118
rect 285784 175596 286364 175624
rect 285784 5166 285812 175596
rect 286704 161474 286732 180118
rect 287060 175636 287112 175642
rect 287060 175578 287112 175584
rect 285876 161446 286732 161474
rect 285876 7614 285904 161446
rect 285864 7608 285916 7614
rect 285864 7550 285916 7556
rect 285772 5160 285824 5166
rect 285772 5102 285824 5108
rect 287072 5030 287100 175578
rect 287164 18630 287192 180118
rect 287704 176996 287756 177002
rect 287704 176938 287756 176944
rect 287716 33794 287744 176938
rect 287808 175642 287836 180118
rect 288452 175658 288480 180118
rect 287796 175636 287848 175642
rect 288452 175630 288572 175658
rect 287796 175578 287848 175584
rect 288440 175568 288492 175574
rect 288440 175510 288492 175516
rect 287704 33788 287756 33794
rect 287704 33730 287756 33736
rect 287152 18624 287204 18630
rect 287152 18566 287204 18572
rect 287060 5024 287112 5030
rect 287060 4966 287112 4972
rect 288452 4962 288480 175510
rect 288544 8090 288572 175630
rect 288636 116618 288664 180118
rect 289280 175574 289308 180118
rect 290200 177546 290228 180118
rect 290292 180118 290674 180146
rect 291028 180118 291134 180146
rect 291304 180118 291686 180146
rect 291764 180118 292238 180146
rect 292698 180118 292804 180146
rect 290188 177540 290240 177546
rect 290188 177482 290240 177488
rect 289268 175568 289320 175574
rect 289268 175510 289320 175516
rect 290292 161474 290320 180118
rect 291028 176730 291056 180118
rect 291200 177404 291252 177410
rect 291200 177346 291252 177352
rect 291016 176724 291068 176730
rect 291016 176666 291068 176672
rect 289832 161446 290320 161474
rect 288624 116612 288676 116618
rect 288624 116554 288676 116560
rect 289832 50386 289860 161446
rect 289820 50380 289872 50386
rect 289820 50322 289872 50328
rect 288992 10464 289044 10470
rect 288992 10406 289044 10412
rect 288532 8084 288584 8090
rect 288532 8026 288584 8032
rect 288440 4956 288492 4962
rect 288440 4898 288492 4904
rect 285692 3454 286640 3482
rect 286612 480 286640 3454
rect 287796 3460 287848 3466
rect 287796 3402 287848 3408
rect 287808 480 287836 3402
rect 289004 480 289032 10406
rect 289820 10396 289872 10402
rect 289820 10338 289872 10344
rect 281878 354 281990 480
rect 281644 326 281990 354
rect 281878 -960 281990 326
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 10338
rect 291212 6914 291240 177346
rect 291304 9178 291332 180118
rect 291764 161474 291792 180118
rect 292580 171828 292632 171834
rect 292580 171770 292632 171776
rect 291396 161446 291792 161474
rect 291396 54534 291424 161446
rect 291384 54528 291436 54534
rect 291384 54470 291436 54476
rect 292592 47734 292620 171770
rect 292776 170406 292804 180118
rect 292868 180118 293250 180146
rect 293328 180118 293710 180146
rect 293972 180118 294262 180146
rect 294340 180118 294814 180146
rect 294892 180118 295274 180146
rect 295352 180118 295826 180146
rect 295904 180118 296286 180146
rect 296732 180118 296838 180146
rect 297390 180118 297496 180146
rect 292764 170400 292816 170406
rect 292764 170342 292816 170348
rect 292868 161474 292896 180118
rect 293328 171834 293356 180118
rect 293316 171828 293368 171834
rect 293316 171770 293368 171776
rect 292776 161446 292896 161474
rect 292776 91798 292804 161446
rect 292764 91792 292816 91798
rect 292764 91734 292816 91740
rect 292580 47728 292632 47734
rect 292580 47670 292632 47676
rect 291292 9172 291344 9178
rect 291292 9114 291344 9120
rect 293684 9036 293736 9042
rect 293684 8978 293736 8984
rect 292580 8968 292632 8974
rect 292580 8910 292632 8916
rect 291212 6886 291424 6914
rect 291396 480 291424 6886
rect 292592 480 292620 8910
rect 293696 480 293724 8978
rect 293972 4894 294000 180118
rect 294340 166994 294368 180118
rect 294064 166966 294368 166994
rect 294064 9110 294092 166966
rect 294892 161474 294920 180118
rect 294156 161446 294920 161474
rect 294156 51746 294184 161446
rect 294144 51740 294196 51746
rect 294144 51682 294196 51688
rect 294144 24132 294196 24138
rect 294144 24074 294196 24080
rect 294156 16574 294184 24074
rect 294156 16546 294920 16574
rect 294052 9104 294104 9110
rect 294052 9046 294104 9052
rect 293960 4888 294012 4894
rect 293960 4830 294012 4836
rect 294892 480 294920 16546
rect 295352 4826 295380 180118
rect 295904 161474 295932 180118
rect 295984 176724 296036 176730
rect 295984 176666 296036 176672
rect 295444 161446 295932 161474
rect 295444 9042 295472 161446
rect 295996 49026 296024 176666
rect 296732 53106 296760 180118
rect 297468 176730 297496 180118
rect 297560 180118 297850 180146
rect 298296 180118 298402 180146
rect 298480 180118 298862 180146
rect 299032 180118 299414 180146
rect 299584 180118 299966 180146
rect 300136 180118 300426 180146
rect 300872 180118 300978 180146
rect 301056 180118 301438 180146
rect 301990 180118 302188 180146
rect 297456 176724 297508 176730
rect 297456 176666 297508 176672
rect 297560 166394 297588 180118
rect 298296 173894 298324 180118
rect 298480 176654 298508 180118
rect 298204 173866 298324 173894
rect 298388 176626 298508 176654
rect 298100 171828 298152 171834
rect 298100 171770 298152 171776
rect 297548 166388 297600 166394
rect 297548 166330 297600 166336
rect 296720 53100 296772 53106
rect 296720 53042 296772 53048
rect 295984 49020 296036 49026
rect 295984 48962 296036 48968
rect 295524 17264 295576 17270
rect 295524 17206 295576 17212
rect 295536 16574 295564 17206
rect 295536 16546 295656 16574
rect 295432 9036 295484 9042
rect 295432 8978 295484 8984
rect 295340 4820 295392 4826
rect 295340 4762 295392 4768
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 297272 13184 297324 13190
rect 297272 13126 297324 13132
rect 297284 480 297312 13126
rect 298112 8974 298140 171770
rect 298204 169130 298232 173866
rect 298204 169102 298324 169130
rect 298192 169040 298244 169046
rect 298192 168982 298244 168988
rect 298204 22846 298232 168982
rect 298296 32434 298324 169102
rect 298388 169046 298416 176626
rect 299032 171834 299060 180118
rect 299020 171828 299072 171834
rect 299020 171770 299072 171776
rect 299480 171828 299532 171834
rect 299480 171770 299532 171776
rect 298376 169040 298428 169046
rect 298376 168982 298428 168988
rect 298284 32428 298336 32434
rect 298284 32370 298336 32376
rect 298284 25560 298336 25566
rect 298284 25502 298336 25508
rect 298192 22840 298244 22846
rect 298192 22782 298244 22788
rect 298100 8968 298152 8974
rect 298100 8910 298152 8916
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298296 354 298324 25502
rect 299492 5098 299520 171770
rect 299584 55894 299612 180118
rect 300032 177540 300084 177546
rect 300032 177482 300084 177488
rect 300044 166994 300072 177482
rect 300136 171834 300164 180118
rect 300872 177546 300900 180118
rect 300860 177540 300912 177546
rect 300860 177482 300912 177488
rect 300124 171828 300176 171834
rect 300124 171770 300176 171776
rect 300044 166966 300164 166994
rect 299572 55888 299624 55894
rect 299572 55830 299624 55836
rect 300136 36582 300164 166966
rect 301056 161474 301084 180118
rect 302160 177410 302188 180118
rect 302252 180118 302542 180146
rect 302712 180118 303002 180146
rect 303264 180118 303554 180146
rect 303632 180118 304014 180146
rect 304092 180118 304566 180146
rect 305012 180118 305118 180146
rect 305288 180118 305578 180146
rect 305840 180118 306130 180146
rect 306392 180118 306590 180146
rect 306668 180118 307142 180146
rect 307588 180118 307694 180146
rect 308154 180118 308260 180146
rect 302148 177404 302200 177410
rect 302148 177346 302200 177352
rect 300872 161446 301084 161474
rect 300872 104174 300900 161446
rect 300860 104168 300912 104174
rect 300860 104110 300912 104116
rect 300124 36576 300176 36582
rect 300124 36518 300176 36524
rect 299572 29640 299624 29646
rect 299572 29582 299624 29588
rect 299480 5092 299532 5098
rect 299480 5034 299532 5040
rect 299584 3534 299612 29582
rect 300860 26920 300912 26926
rect 300860 26862 300912 26868
rect 299664 22772 299716 22778
rect 299664 22714 299716 22720
rect 299572 3528 299624 3534
rect 299572 3470 299624 3476
rect 299676 480 299704 22714
rect 300872 16574 300900 26862
rect 300872 16546 301544 16574
rect 300768 3528 300820 3534
rect 300768 3470 300820 3476
rect 300780 480 300808 3470
rect 298438 354 298550 480
rect 298296 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16546
rect 302252 9382 302280 180118
rect 302332 175636 302384 175642
rect 302332 175578 302384 175584
rect 302344 24138 302372 175578
rect 302712 161474 302740 180118
rect 303264 175642 303292 180118
rect 303252 175636 303304 175642
rect 303252 175578 303304 175584
rect 302436 161446 302740 161474
rect 302436 57254 302464 161446
rect 302424 57248 302476 57254
rect 302424 57190 302476 57196
rect 303632 42226 303660 180118
rect 304092 161474 304120 180118
rect 304264 176724 304316 176730
rect 304264 176666 304316 176672
rect 303724 161446 304120 161474
rect 303724 60042 303752 161446
rect 303712 60036 303764 60042
rect 303712 59978 303764 59984
rect 303620 42220 303672 42226
rect 303620 42162 303672 42168
rect 302332 24132 302384 24138
rect 302332 24074 302384 24080
rect 304276 17338 304304 176666
rect 305012 25566 305040 180118
rect 305184 175636 305236 175642
rect 305184 175578 305236 175584
rect 305196 58682 305224 175578
rect 305288 129062 305316 180118
rect 305840 175642 305868 180118
rect 305828 175636 305880 175642
rect 305828 175578 305880 175584
rect 305276 129056 305328 129062
rect 305276 128998 305328 129004
rect 305184 58676 305236 58682
rect 305184 58618 305236 58624
rect 305092 31068 305144 31074
rect 305092 31010 305144 31016
rect 305000 25560 305052 25566
rect 305000 25502 305052 25508
rect 304264 17332 304316 17338
rect 304264 17274 304316 17280
rect 305104 16574 305132 31010
rect 306392 26994 306420 180118
rect 306668 161474 306696 180118
rect 307024 177472 307076 177478
rect 307024 177414 307076 177420
rect 306484 161446 306696 161474
rect 306484 152522 306512 161446
rect 306472 152516 306524 152522
rect 306472 152458 306524 152464
rect 306380 26988 306432 26994
rect 306380 26930 306432 26936
rect 305104 16546 305592 16574
rect 303160 13116 303212 13122
rect 303160 13058 303212 13064
rect 302240 9376 302292 9382
rect 302240 9318 302292 9324
rect 303172 480 303200 13058
rect 304356 6248 304408 6254
rect 304356 6190 304408 6196
rect 304368 480 304396 6190
rect 305564 480 305592 16546
rect 306380 14544 306432 14550
rect 306380 14486 306432 14492
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 354 306420 14486
rect 307036 13122 307064 177414
rect 307588 176730 307616 180118
rect 308232 177818 308260 180118
rect 308324 180118 308706 180146
rect 309166 180118 309272 180146
rect 308220 177812 308272 177818
rect 308220 177754 308272 177760
rect 307576 176724 307628 176730
rect 307576 176666 307628 176672
rect 308324 163606 308352 180118
rect 309244 175658 309272 180118
rect 309612 180118 309718 180146
rect 309796 180118 310270 180146
rect 310624 180118 310730 180146
rect 310808 180118 311282 180146
rect 311360 180118 311742 180146
rect 312004 180118 312294 180146
rect 312464 180118 312846 180146
rect 313306 180118 313412 180146
rect 309612 176050 309640 180118
rect 309600 176044 309652 176050
rect 309600 175986 309652 175992
rect 309152 175630 309272 175658
rect 308312 163600 308364 163606
rect 308312 163542 308364 163548
rect 309152 61402 309180 175630
rect 309796 174706 309824 180118
rect 309968 177540 310020 177546
rect 309968 177482 310020 177488
rect 309876 176724 309928 176730
rect 309876 176666 309928 176672
rect 309244 174678 309824 174706
rect 309244 153950 309272 174678
rect 309888 174570 309916 176666
rect 309796 174542 309916 174570
rect 309232 153944 309284 153950
rect 309232 153886 309284 153892
rect 309140 61396 309192 61402
rect 309140 61338 309192 61344
rect 307760 35216 307812 35222
rect 307760 35158 307812 35164
rect 307024 13116 307076 13122
rect 307024 13058 307076 13064
rect 307772 3534 307800 35158
rect 307852 21480 307904 21486
rect 307852 21422 307904 21428
rect 307864 16574 307892 21422
rect 307864 16546 307984 16574
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 307956 480 307984 16546
rect 309692 15972 309744 15978
rect 309692 15914 309744 15920
rect 309704 6914 309732 15914
rect 309796 14550 309824 174542
rect 309980 161474 310008 177482
rect 310520 175636 310572 175642
rect 310520 175578 310572 175584
rect 309888 161446 310008 161474
rect 309888 44878 309916 161446
rect 309876 44872 309928 44878
rect 309876 44814 309928 44820
rect 309784 14544 309836 14550
rect 309784 14486 309836 14492
rect 310532 10742 310560 175578
rect 310624 19990 310652 180118
rect 310808 149802 310836 180118
rect 311360 175642 311388 180118
rect 311348 175636 311400 175642
rect 311348 175578 311400 175584
rect 311900 175636 311952 175642
rect 311900 175578 311952 175584
rect 310796 149796 310848 149802
rect 310796 149738 310848 149744
rect 310704 32496 310756 32502
rect 310704 32438 310756 32444
rect 310612 19984 310664 19990
rect 310612 19926 310664 19932
rect 310716 16574 310744 32438
rect 310716 16546 311480 16574
rect 310520 10736 310572 10742
rect 310520 10678 310572 10684
rect 309704 6886 309824 6914
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 306718 354 306830 480
rect 306392 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 311452 480 311480 16546
rect 311912 6458 311940 175578
rect 312004 164966 312032 180118
rect 312464 175642 312492 180118
rect 312544 177404 312596 177410
rect 312544 177346 312596 177352
rect 312452 175636 312504 175642
rect 312452 175578 312504 175584
rect 311992 164960 312044 164966
rect 311992 164902 312044 164908
rect 312556 127634 312584 177346
rect 313384 175658 313412 180118
rect 313292 175630 313412 175658
rect 313476 180118 313858 180146
rect 313936 180118 314318 180146
rect 314764 180118 314870 180146
rect 314948 180118 315422 180146
rect 315882 180118 315988 180146
rect 312544 127628 312596 127634
rect 312544 127570 312596 127576
rect 311992 37936 312044 37942
rect 311992 37878 312044 37884
rect 312004 16574 312032 37878
rect 312004 16546 312216 16574
rect 311900 6452 311952 6458
rect 311900 6394 311952 6400
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313292 10674 313320 175630
rect 313372 175568 313424 175574
rect 313372 175510 313424 175516
rect 313280 10668 313332 10674
rect 313280 10610 313332 10616
rect 313384 6390 313412 175510
rect 313476 155310 313504 180118
rect 313936 175574 313964 180118
rect 313924 175568 313976 175574
rect 313924 175510 313976 175516
rect 314764 171902 314792 180118
rect 314752 171896 314804 171902
rect 314752 171838 314804 171844
rect 314948 161474 314976 180118
rect 315960 177410 315988 180118
rect 316144 180118 316434 180146
rect 316512 180118 316894 180146
rect 317446 180118 317552 180146
rect 315948 177404 316000 177410
rect 315948 177346 316000 177352
rect 316040 175976 316092 175982
rect 316040 175918 316092 175924
rect 314672 161446 314976 161474
rect 314672 156738 314700 161446
rect 314660 156732 314712 156738
rect 314660 156674 314712 156680
rect 313464 155304 313516 155310
rect 313464 155246 313516 155252
rect 313832 11824 313884 11830
rect 313832 11766 313884 11772
rect 313372 6384 313424 6390
rect 313372 6326 313424 6332
rect 313844 480 313872 11766
rect 314660 10328 314712 10334
rect 314660 10270 314712 10276
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 10270
rect 316052 3534 316080 175918
rect 316144 10606 316172 180118
rect 316512 161474 316540 180118
rect 317524 175658 317552 180118
rect 316236 161446 316540 161474
rect 317432 175630 317552 175658
rect 317616 180118 317998 180146
rect 318168 180118 318458 180146
rect 318904 180118 319010 180146
rect 319088 180118 319470 180146
rect 320022 180118 320128 180146
rect 316236 160818 316264 161446
rect 316224 160812 316276 160818
rect 316224 160754 316276 160760
rect 316224 14476 316276 14482
rect 316224 14418 316276 14424
rect 316132 10600 316184 10606
rect 316132 10542 316184 10548
rect 316040 3528 316092 3534
rect 316040 3470 316092 3476
rect 316236 480 316264 14418
rect 317432 6322 317460 175630
rect 317512 175568 317564 175574
rect 317512 175510 317564 175516
rect 317420 6316 317472 6322
rect 317420 6258 317472 6264
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 317340 480 317368 3470
rect 317524 3262 317552 175510
rect 317616 10538 317644 180118
rect 318168 175574 318196 180118
rect 318904 176730 318932 180118
rect 318892 176724 318944 176730
rect 318892 176666 318944 176672
rect 318156 175568 318208 175574
rect 318156 175510 318208 175516
rect 319088 162246 319116 180118
rect 320100 177750 320128 180118
rect 320192 180118 320574 180146
rect 320652 180118 321034 180146
rect 321586 180118 321692 180146
rect 320088 177744 320140 177750
rect 320088 177686 320140 177692
rect 319076 162240 319128 162246
rect 319076 162182 319128 162188
rect 318800 39364 318852 39370
rect 318800 39306 318852 39312
rect 318812 16574 318840 39306
rect 318812 16546 319760 16574
rect 317604 10532 317656 10538
rect 317604 10474 317656 10480
rect 318524 6588 318576 6594
rect 318524 6530 318576 6536
rect 317512 3256 317564 3262
rect 317512 3198 317564 3204
rect 318536 480 318564 6530
rect 319732 480 319760 16546
rect 320192 6254 320220 180118
rect 320652 161474 320680 180118
rect 320824 177404 320876 177410
rect 320824 177346 320876 177352
rect 320284 161446 320680 161474
rect 320284 10470 320312 161446
rect 320836 43450 320864 177346
rect 321664 176654 321692 180118
rect 321572 176626 321692 176654
rect 321756 180118 322046 180146
rect 322216 180118 322598 180146
rect 323150 180118 323256 180146
rect 320824 43444 320876 43450
rect 320824 43386 320876 43392
rect 320364 18692 320416 18698
rect 320364 18634 320416 18640
rect 320376 16574 320404 18634
rect 320376 16546 320496 16574
rect 320272 10464 320324 10470
rect 320272 10406 320324 10412
rect 320180 6248 320232 6254
rect 320180 6190 320232 6196
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 321572 3330 321600 176626
rect 321652 171148 321704 171154
rect 321652 171090 321704 171096
rect 321664 10402 321692 171090
rect 321756 148442 321784 180118
rect 322216 171154 322244 180118
rect 323228 177682 323256 180118
rect 323320 180118 323610 180146
rect 323872 180118 324162 180146
rect 324332 180118 324622 180146
rect 324700 180118 325174 180146
rect 325726 180118 325832 180146
rect 326186 180118 326568 180146
rect 326738 180118 327028 180146
rect 327290 180118 327396 180146
rect 323216 177676 323268 177682
rect 323216 177618 323268 177624
rect 322940 171828 322992 171834
rect 322940 171770 322992 171776
rect 322204 171148 322256 171154
rect 322204 171090 322256 171096
rect 321744 148436 321796 148442
rect 321744 148378 321796 148384
rect 321652 10396 321704 10402
rect 321652 10338 321704 10344
rect 322952 10334 322980 171770
rect 323320 161474 323348 180118
rect 323584 176724 323636 176730
rect 323584 176666 323636 176672
rect 323044 161446 323348 161474
rect 323044 35222 323072 161446
rect 323124 40724 323176 40730
rect 323124 40666 323176 40672
rect 323032 35216 323084 35222
rect 323032 35158 323084 35164
rect 322940 10328 322992 10334
rect 322940 10270 322992 10276
rect 322112 6520 322164 6526
rect 322112 6462 322164 6468
rect 321560 3324 321612 3330
rect 321560 3266 321612 3272
rect 322124 480 322152 6462
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 323136 354 323164 40666
rect 323596 29646 323624 176666
rect 323872 171834 323900 180118
rect 323860 171828 323912 171834
rect 323860 171770 323912 171776
rect 323584 29640 323636 29646
rect 323584 29582 323636 29588
rect 324332 3398 324360 180118
rect 324412 173188 324464 173194
rect 324412 173130 324464 173136
rect 324424 3602 324452 173130
rect 324700 161474 324728 180118
rect 325804 161474 325832 180118
rect 326540 177614 326568 180118
rect 326528 177608 326580 177614
rect 326528 177550 326580 177556
rect 327000 176730 327028 180118
rect 326988 176724 327040 176730
rect 326988 176666 327040 176672
rect 327368 176662 327396 180118
rect 327460 180118 327750 180146
rect 327920 180118 328302 180146
rect 328472 180118 328762 180146
rect 329314 180118 329696 180146
rect 329866 180118 329972 180146
rect 327356 176656 327408 176662
rect 327356 176598 327408 176604
rect 327460 172122 327488 180118
rect 327540 176656 327592 176662
rect 327540 176598 327592 176604
rect 324516 161446 324728 161474
rect 325712 161446 325832 161474
rect 327092 172094 327488 172122
rect 324516 147014 324544 161446
rect 324504 147008 324556 147014
rect 324504 146950 324556 146956
rect 325712 124914 325740 161446
rect 325700 124908 325752 124914
rect 325700 124850 325752 124856
rect 325700 46232 325752 46238
rect 325700 46174 325752 46180
rect 324504 28280 324556 28286
rect 324504 28222 324556 28228
rect 324412 3596 324464 3602
rect 324412 3538 324464 3544
rect 324516 3482 324544 28222
rect 325712 16574 325740 46174
rect 325712 16546 326384 16574
rect 325608 3596 325660 3602
rect 325608 3538 325660 3544
rect 324424 3454 324544 3482
rect 324320 3392 324372 3398
rect 324320 3334 324372 3340
rect 324424 480 324452 3454
rect 325620 480 325648 3538
rect 323278 354 323390 480
rect 323136 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 327092 4146 327120 172094
rect 327172 171828 327224 171834
rect 327172 171770 327224 171776
rect 327184 93158 327212 171770
rect 327552 161474 327580 176598
rect 327920 171834 327948 180118
rect 327908 171828 327960 171834
rect 327908 171770 327960 171776
rect 327276 161446 327580 161474
rect 327276 158098 327304 161446
rect 328472 159458 328500 180118
rect 329668 177546 329696 180118
rect 329656 177540 329708 177546
rect 329656 177482 329708 177488
rect 329104 177336 329156 177342
rect 329104 177278 329156 177284
rect 328460 159452 328512 159458
rect 328460 159394 328512 159400
rect 327264 158092 327316 158098
rect 327264 158034 327316 158040
rect 327172 93152 327224 93158
rect 327172 93094 327224 93100
rect 327172 20052 327224 20058
rect 327172 19994 327224 20000
rect 327184 16574 327212 19994
rect 327184 16546 328040 16574
rect 327080 4140 327132 4146
rect 327080 4082 327132 4088
rect 328012 480 328040 16546
rect 329116 11762 329144 177278
rect 329196 176724 329248 176730
rect 329196 176666 329248 176672
rect 329208 31074 329236 176666
rect 329944 176654 329972 180118
rect 329852 176626 329972 176654
rect 330036 180118 330326 180146
rect 330496 180118 330878 180146
rect 331232 180118 331338 180146
rect 331416 180118 331890 180146
rect 332442 180118 332548 180146
rect 332902 180118 333192 180146
rect 329852 145586 329880 176626
rect 329932 171148 329984 171154
rect 329932 171090 329984 171096
rect 329840 145580 329892 145586
rect 329840 145522 329892 145528
rect 329840 123480 329892 123486
rect 329840 123422 329892 123428
rect 329196 31068 329248 31074
rect 329196 31010 329248 31016
rect 329104 11756 329156 11762
rect 329104 11698 329156 11704
rect 329196 6180 329248 6186
rect 329196 6122 329248 6128
rect 329208 480 329236 6122
rect 329852 3482 329880 123422
rect 329944 4078 329972 171090
rect 330036 123486 330064 180118
rect 330496 171154 330524 180118
rect 330484 171148 330536 171154
rect 330484 171090 330536 171096
rect 330024 123480 330076 123486
rect 330024 123422 330076 123428
rect 331232 28286 331260 180118
rect 331416 122126 331444 180118
rect 332520 177478 332548 180118
rect 332508 177472 332560 177478
rect 332508 177414 332560 177420
rect 333164 177138 333192 180118
rect 333348 180118 333454 180146
rect 333532 180118 333914 180146
rect 334084 180118 334466 180146
rect 334636 180118 335018 180146
rect 335372 180118 335478 180146
rect 335556 180118 336030 180146
rect 336108 180118 336490 180146
rect 336752 180118 337042 180146
rect 337488 180118 337594 180146
rect 337672 180118 338054 180146
rect 338500 180118 338606 180146
rect 338684 180118 339066 180146
rect 339512 180118 339618 180146
rect 339880 180118 340170 180146
rect 340248 180118 340630 180146
rect 341076 180118 341182 180146
rect 341352 180118 341642 180146
rect 341904 180118 342194 180146
rect 342364 180118 342746 180146
rect 342824 180118 343206 180146
rect 343652 180118 343758 180146
rect 343836 180118 344218 180146
rect 344480 180118 344770 180146
rect 345124 180118 345322 180146
rect 345400 180118 345782 180146
rect 345952 180118 346334 180146
rect 346504 180118 346794 180146
rect 347056 180118 347346 180146
rect 347898 180118 348004 180146
rect 348358 180118 348464 180146
rect 333152 177132 333204 177138
rect 333152 177074 333204 177080
rect 333348 173262 333376 180118
rect 333336 173256 333388 173262
rect 333336 173198 333388 173204
rect 333532 161474 333560 180118
rect 333980 174548 334032 174554
rect 333980 174490 334032 174496
rect 332612 161446 333560 161474
rect 331404 122120 331456 122126
rect 331404 122062 331456 122068
rect 331220 28280 331272 28286
rect 331220 28222 331272 28228
rect 331220 11756 331272 11762
rect 331220 11698 331272 11704
rect 329932 4072 329984 4078
rect 329932 4014 329984 4020
rect 329852 3454 330432 3482
rect 330404 480 330432 3454
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 11698
rect 332612 4010 332640 161446
rect 333992 16574 334020 174490
rect 334084 94518 334112 180118
rect 334636 161474 334664 180118
rect 335372 177410 335400 180118
rect 335360 177404 335412 177410
rect 335360 177346 335412 177352
rect 335556 175794 335584 180118
rect 334176 161446 334664 161474
rect 335372 175766 335584 175794
rect 334176 120766 334204 161446
rect 334164 120760 334216 120766
rect 334164 120702 334216 120708
rect 334072 94512 334124 94518
rect 334072 94454 334124 94460
rect 333992 16546 334664 16574
rect 332692 15904 332744 15910
rect 332692 15846 332744 15852
rect 332600 4004 332652 4010
rect 332600 3946 332652 3952
rect 332704 3602 332732 15846
rect 332784 11688 332836 11694
rect 332784 11630 332836 11636
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 332796 3482 332824 11630
rect 333888 3596 333940 3602
rect 333888 3538 333940 3544
rect 332704 3454 332824 3482
rect 332704 480 332732 3454
rect 333900 480 333928 3538
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 16546
rect 335372 8022 335400 175766
rect 336108 175658 336136 180118
rect 336188 177132 336240 177138
rect 336188 177074 336240 177080
rect 335556 175630 336136 175658
rect 335556 46238 335584 175630
rect 336200 161474 336228 177074
rect 336016 161446 336228 161474
rect 336016 144226 336044 161446
rect 336004 144220 336056 144226
rect 336004 144162 336056 144168
rect 335544 46232 335596 46238
rect 335544 46174 335596 46180
rect 335452 33788 335504 33794
rect 335452 33730 335504 33736
rect 335464 16574 335492 33730
rect 335464 16546 336320 16574
rect 335360 8016 335412 8022
rect 335360 7958 335412 7964
rect 336292 480 336320 16546
rect 336752 3942 336780 180118
rect 337488 176730 337516 180118
rect 337476 176724 337528 176730
rect 337476 176666 337528 176672
rect 337672 169114 337700 180118
rect 338500 177342 338528 180118
rect 338488 177336 338540 177342
rect 338488 177278 338540 177284
rect 337660 169108 337712 169114
rect 337660 169050 337712 169056
rect 338684 161474 338712 180118
rect 338764 177812 338816 177818
rect 338764 177754 338816 177760
rect 338132 161446 338712 161474
rect 336832 21412 336884 21418
rect 336832 21354 336884 21360
rect 336844 16574 336872 21354
rect 336844 16546 337056 16574
rect 336740 3936 336792 3942
rect 336740 3878 336792 3884
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338132 7954 338160 161446
rect 338776 18698 338804 177754
rect 338856 176724 338908 176730
rect 338856 176666 338908 176672
rect 338868 142866 338896 176666
rect 339512 175624 339540 180118
rect 339512 175596 339632 175624
rect 339500 175500 339552 175506
rect 339500 175442 339552 175448
rect 338856 142860 338908 142866
rect 338856 142802 338908 142808
rect 338764 18692 338816 18698
rect 338764 18634 338816 18640
rect 338120 7948 338172 7954
rect 338120 7890 338172 7896
rect 338672 5228 338724 5234
rect 338672 5170 338724 5176
rect 338684 480 338712 5170
rect 339512 3874 339540 175442
rect 339604 119406 339632 175596
rect 339880 175506 339908 180118
rect 339868 175500 339920 175506
rect 339868 175442 339920 175448
rect 340248 161474 340276 180118
rect 340972 175704 341024 175710
rect 340972 175646 341024 175652
rect 340880 175636 340932 175642
rect 340880 175578 340932 175584
rect 339696 161446 340276 161474
rect 339592 119400 339644 119406
rect 339592 119342 339644 119348
rect 339696 7886 339724 161446
rect 339684 7880 339736 7886
rect 339684 7822 339736 7828
rect 339868 7676 339920 7682
rect 339868 7618 339920 7624
rect 339500 3868 339552 3874
rect 339500 3810 339552 3816
rect 339880 480 339908 7618
rect 340892 3806 340920 175578
rect 340984 13258 341012 175646
rect 340972 13252 341024 13258
rect 340972 13194 341024 13200
rect 340972 13116 341024 13122
rect 340972 13058 341024 13064
rect 340880 3800 340932 3806
rect 340880 3742 340932 3748
rect 340984 480 341012 13058
rect 341076 12102 341104 180118
rect 341352 175642 341380 180118
rect 341904 175710 341932 180118
rect 341892 175704 341944 175710
rect 341892 175646 341944 175652
rect 341340 175636 341392 175642
rect 341340 175578 341392 175584
rect 342260 175636 342312 175642
rect 342260 175578 342312 175584
rect 341156 13252 341208 13258
rect 341156 13194 341208 13200
rect 341064 12096 341116 12102
rect 341064 12038 341116 12044
rect 341168 7818 341196 13194
rect 341156 7812 341208 7818
rect 341156 7754 341208 7760
rect 342168 5160 342220 5166
rect 342168 5102 342220 5108
rect 342180 480 342208 5102
rect 342272 3738 342300 175578
rect 342364 12034 342392 180118
rect 342824 175642 342852 180118
rect 343652 177206 343680 180118
rect 343640 177200 343692 177206
rect 343640 177142 343692 177148
rect 342812 175636 342864 175642
rect 342812 175578 342864 175584
rect 343640 175636 343692 175642
rect 343640 175578 343692 175584
rect 342352 12028 342404 12034
rect 342352 11970 342404 11976
rect 343364 7608 343416 7614
rect 343364 7550 343416 7556
rect 342260 3732 342312 3738
rect 342260 3674 342312 3680
rect 343376 480 343404 7550
rect 343652 3670 343680 175578
rect 343836 117978 343864 180118
rect 344480 175642 344508 180118
rect 344468 175636 344520 175642
rect 344468 175578 344520 175584
rect 345020 175636 345072 175642
rect 345020 175578 345072 175584
rect 343824 117972 343876 117978
rect 343824 117914 343876 117920
rect 343732 18624 343784 18630
rect 343732 18566 343784 18572
rect 343744 16574 343772 18566
rect 343744 16546 344600 16574
rect 343640 3664 343692 3670
rect 343640 3606 343692 3612
rect 344572 480 344600 16546
rect 345032 3534 345060 175578
rect 345124 7750 345152 180118
rect 345400 161474 345428 180118
rect 345952 175642 345980 180118
rect 345940 175636 345992 175642
rect 345940 175578 345992 175584
rect 346400 173868 346452 173874
rect 346400 173810 346452 173816
rect 345216 161446 345428 161474
rect 345216 11966 345244 161446
rect 345204 11960 345256 11966
rect 345204 11902 345256 11908
rect 345112 7744 345164 7750
rect 345112 7686 345164 7692
rect 346412 7682 346440 173810
rect 346504 14482 346532 180118
rect 346952 177200 347004 177206
rect 346952 177142 347004 177148
rect 346964 171134 346992 177142
rect 347056 173874 347084 180118
rect 347780 175636 347832 175642
rect 347780 175578 347832 175584
rect 347044 173868 347096 173874
rect 347044 173810 347096 173816
rect 346964 171106 347084 171134
rect 347056 33794 347084 171106
rect 347792 141438 347820 175578
rect 347976 161474 348004 180118
rect 348436 174622 348464 180118
rect 348528 180118 348910 180146
rect 349264 180118 349370 180146
rect 349448 180118 349922 180146
rect 350184 180118 350474 180146
rect 350552 180118 350934 180146
rect 351486 180118 351776 180146
rect 351946 180118 352052 180146
rect 348528 175642 348556 180118
rect 348516 175636 348568 175642
rect 348516 175578 348568 175584
rect 349160 175636 349212 175642
rect 349160 175578 349212 175584
rect 348424 174616 348476 174622
rect 348424 174558 348476 174564
rect 347884 161446 348004 161474
rect 347780 141432 347832 141438
rect 347780 141374 347832 141380
rect 347884 116686 347912 161446
rect 347872 116680 347924 116686
rect 347872 116622 347924 116628
rect 347780 116612 347832 116618
rect 347780 116554 347832 116560
rect 347044 33788 347096 33794
rect 347044 33730 347096 33736
rect 347792 16574 347820 116554
rect 347792 16546 348096 16574
rect 346492 14476 346544 14482
rect 346492 14418 346544 14424
rect 346952 8084 347004 8090
rect 346952 8026 347004 8032
rect 346400 7676 346452 7682
rect 346400 7618 346452 7624
rect 345756 5024 345808 5030
rect 345756 4966 345808 4972
rect 345020 3528 345072 3534
rect 345020 3470 345072 3476
rect 345768 480 345796 4966
rect 346964 480 346992 8026
rect 348068 480 348096 16546
rect 349172 7614 349200 175578
rect 349264 11898 349292 180118
rect 349344 36576 349396 36582
rect 349344 36518 349396 36524
rect 349252 11892 349304 11898
rect 349252 11834 349304 11840
rect 349160 7608 349212 7614
rect 349160 7550 349212 7556
rect 349356 6914 349384 36518
rect 349448 15910 349476 180118
rect 350184 175642 350212 180118
rect 350172 175636 350224 175642
rect 350172 175578 350224 175584
rect 350552 115258 350580 180118
rect 351748 173194 351776 180118
rect 351736 173188 351788 173194
rect 351736 173130 351788 173136
rect 352024 166994 352052 180118
rect 351932 166966 352052 166994
rect 352116 180118 352498 180146
rect 353050 180118 353248 180146
rect 353510 180118 353616 180146
rect 350540 115252 350592 115258
rect 350540 115194 350592 115200
rect 350540 50380 350592 50386
rect 350540 50322 350592 50328
rect 350552 16574 350580 50322
rect 351932 36582 351960 166966
rect 352116 161474 352144 180118
rect 353220 171698 353248 180118
rect 353300 171828 353352 171834
rect 353300 171770 353352 171776
rect 353208 171692 353260 171698
rect 353208 171634 353260 171640
rect 352024 161446 352144 161474
rect 351920 36576 351972 36582
rect 351920 36518 351972 36524
rect 350552 16546 351224 16574
rect 349436 15904 349488 15910
rect 349436 15846 349488 15852
rect 349356 6886 350488 6914
rect 349252 4956 349304 4962
rect 349252 4898 349304 4904
rect 349264 480 349292 4898
rect 350460 480 350488 6886
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351196 354 351224 16546
rect 352024 11830 352052 161446
rect 352104 49020 352156 49026
rect 352104 48962 352156 48968
rect 352116 16574 352144 48962
rect 352116 16546 352880 16574
rect 352012 11824 352064 11830
rect 352012 11766 352064 11772
rect 352852 480 352880 16546
rect 353312 11762 353340 171770
rect 353392 171760 353444 171766
rect 353392 171702 353444 171708
rect 353404 21418 353432 171702
rect 353588 161474 353616 180118
rect 353680 180118 354062 180146
rect 354232 180118 354522 180146
rect 354968 180118 355074 180146
rect 355152 180118 355626 180146
rect 353680 171834 353708 180118
rect 353668 171828 353720 171834
rect 353668 171770 353720 171776
rect 354232 171766 354260 180118
rect 354968 176730 354996 180118
rect 354956 176724 355008 176730
rect 354956 176666 355008 176672
rect 354220 171760 354272 171766
rect 354220 171702 354272 171708
rect 355152 161474 355180 180118
rect 356152 171828 356204 171834
rect 356152 171770 356204 171776
rect 356060 170400 356112 170406
rect 356060 170342 356112 170348
rect 353496 161446 353616 161474
rect 354692 161446 355180 161474
rect 353496 140078 353524 161446
rect 353484 140072 353536 140078
rect 353484 140014 353536 140020
rect 354692 113830 354720 161446
rect 354680 113824 354732 113830
rect 354680 113766 354732 113772
rect 354680 54528 354732 54534
rect 354680 54470 354732 54476
rect 353392 21412 353444 21418
rect 353392 21354 353444 21360
rect 354692 16574 354720 54470
rect 354692 16546 355272 16574
rect 353300 11756 353352 11762
rect 353300 11698 353352 11704
rect 354036 9172 354088 9178
rect 354036 9114 354088 9120
rect 354048 480 354076 9114
rect 355244 480 355272 16546
rect 356072 6914 356100 170342
rect 356164 13326 356192 171770
rect 356348 170406 356376 180254
rect 356440 180118 356638 180146
rect 356808 180118 357098 180146
rect 357650 180118 357756 180146
rect 356336 170400 356388 170406
rect 356336 170342 356388 170348
rect 356440 166994 356468 180118
rect 356808 171834 356836 180118
rect 357728 176662 357756 180118
rect 357820 180118 358202 180146
rect 358280 180118 358662 180146
rect 358924 180118 359214 180146
rect 359384 180118 359766 180146
rect 360226 180118 360332 180146
rect 357716 176656 357768 176662
rect 357716 176598 357768 176604
rect 356796 171828 356848 171834
rect 356796 171770 356848 171776
rect 357440 171828 357492 171834
rect 357440 171770 357492 171776
rect 356256 166966 356468 166994
rect 356256 137290 356284 166966
rect 356244 137284 356296 137290
rect 356244 137226 356296 137232
rect 357452 47598 357480 171770
rect 357820 166994 357848 180118
rect 357900 176656 357952 176662
rect 357900 176598 357952 176604
rect 357544 166966 357848 166994
rect 357544 135930 357572 166966
rect 357912 161474 357940 176598
rect 358280 171834 358308 180118
rect 358268 171828 358320 171834
rect 358268 171770 358320 171776
rect 358924 169046 358952 180118
rect 358912 169040 358964 169046
rect 358912 168982 358964 168988
rect 359384 166994 359412 180118
rect 359464 176724 359516 176730
rect 359464 176666 359516 176672
rect 357636 161446 357940 161474
rect 358832 166966 359412 166994
rect 357532 135924 357584 135930
rect 357532 135866 357584 135872
rect 357636 91798 357664 161446
rect 357532 91792 357584 91798
rect 357532 91734 357584 91740
rect 357624 91792 357676 91798
rect 357624 91734 357676 91740
rect 357440 47592 357492 47598
rect 357440 47534 357492 47540
rect 356152 13320 356204 13326
rect 356152 13262 356204 13268
rect 356072 6886 356376 6914
rect 356348 480 356376 6886
rect 357544 480 357572 91734
rect 357624 47728 357676 47734
rect 357624 47670 357676 47676
rect 357636 16574 357664 47670
rect 358832 37942 358860 166966
rect 358820 37936 358872 37942
rect 358820 37878 358872 37884
rect 359476 22778 359504 176666
rect 360304 174434 360332 180118
rect 360212 174406 360332 174434
rect 360396 180118 360778 180146
rect 360856 180118 361238 180146
rect 361592 180118 361790 180146
rect 361868 180118 362342 180146
rect 362802 180118 362908 180146
rect 359464 22772 359516 22778
rect 359464 22714 359516 22720
rect 357636 16546 358768 16574
rect 358740 480 358768 16546
rect 360212 13258 360240 174406
rect 360396 174298 360424 180118
rect 360304 174270 360424 174298
rect 360200 13252 360252 13258
rect 360200 13194 360252 13200
rect 360304 5030 360332 174270
rect 360856 161474 360884 180118
rect 360396 161446 360884 161474
rect 360396 134570 360424 161446
rect 360384 134564 360436 134570
rect 360384 134506 360436 134512
rect 361592 111110 361620 180118
rect 361868 167686 361896 180118
rect 362880 176730 362908 180118
rect 363064 180118 363354 180146
rect 363432 180118 363814 180146
rect 364366 180118 364472 180146
rect 362868 176724 362920 176730
rect 362868 176666 362920 176672
rect 362960 175636 363012 175642
rect 362960 175578 363012 175584
rect 361856 167680 361908 167686
rect 361856 167622 361908 167628
rect 361580 111104 361632 111110
rect 361580 111046 361632 111052
rect 361580 51740 361632 51746
rect 361580 51682 361632 51688
rect 361592 16574 361620 51682
rect 361592 16546 361896 16574
rect 361120 9104 361172 9110
rect 361120 9046 361172 9052
rect 360292 5024 360344 5030
rect 360292 4966 360344 4972
rect 359924 4888 359976 4894
rect 359924 4830 359976 4836
rect 359936 480 359964 4830
rect 361132 480 361160 9046
rect 351614 354 351726 480
rect 351196 326 351726 354
rect 351614 -960 351726 326
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 361868 354 361896 16546
rect 362972 4962 363000 175578
rect 363064 13190 363092 180118
rect 363432 175642 363460 180118
rect 363604 176724 363656 176730
rect 363604 176666 363656 176672
rect 363420 175636 363472 175642
rect 363420 175578 363472 175584
rect 363616 133210 363644 176666
rect 364444 175658 364472 180118
rect 364352 175630 364472 175658
rect 364536 180118 364918 180146
rect 364996 180118 365378 180146
rect 365732 180118 365930 180146
rect 366008 180118 366390 180146
rect 366468 180118 366942 180146
rect 367112 180118 367494 180146
rect 367572 180118 367954 180146
rect 368506 180118 368612 180146
rect 363604 133204 363656 133210
rect 363604 133146 363656 133152
rect 364352 131782 364380 175630
rect 364536 174434 364564 180118
rect 364444 174406 364564 174434
rect 364340 131776 364392 131782
rect 364340 131718 364392 131724
rect 363052 13184 363104 13190
rect 363052 13126 363104 13132
rect 364444 13122 364472 174406
rect 364996 161474 365024 180118
rect 364536 161446 365024 161474
rect 364536 17270 364564 161446
rect 365732 39370 365760 180118
rect 366008 175658 366036 180118
rect 365824 175630 366036 175658
rect 365824 109750 365852 175630
rect 366468 166326 366496 180118
rect 366456 166320 366508 166326
rect 366456 166262 366508 166268
rect 365812 109744 365864 109750
rect 365812 109686 365864 109692
rect 365812 53100 365864 53106
rect 365812 53042 365864 53048
rect 365720 39364 365772 39370
rect 365720 39306 365772 39312
rect 365720 17332 365772 17338
rect 365720 17274 365772 17280
rect 364524 17264 364576 17270
rect 364524 17206 364576 17212
rect 364432 13116 364484 13122
rect 364432 13058 364484 13064
rect 364616 9036 364668 9042
rect 364616 8978 364668 8984
rect 362960 4956 363012 4962
rect 362960 4898 363012 4904
rect 363512 4820 363564 4826
rect 363512 4762 363564 4768
rect 363524 480 363552 4762
rect 364628 480 364656 8978
rect 365732 3466 365760 17274
rect 365720 3460 365772 3466
rect 365720 3402 365772 3408
rect 365824 480 365852 53042
rect 367112 9314 367140 180118
rect 367192 166388 367244 166394
rect 367192 166330 367244 166336
rect 367204 16574 367232 166330
rect 367572 161474 367600 180118
rect 368584 174570 368612 180118
rect 368860 180118 368966 180146
rect 369044 180118 369518 180146
rect 369872 180118 370070 180146
rect 370148 180118 370530 180146
rect 370700 180118 371082 180146
rect 371252 180118 371542 180146
rect 371620 180118 372094 180146
rect 372646 180118 372752 180146
rect 368860 176730 368888 180118
rect 368848 176724 368900 176730
rect 368848 176666 368900 176672
rect 368492 174542 368612 174570
rect 368492 164898 368520 174542
rect 368480 164892 368532 164898
rect 368480 164834 368532 164840
rect 369044 161474 369072 180118
rect 367296 161446 367600 161474
rect 368584 161446 369072 161474
rect 367296 146946 367324 161446
rect 367284 146940 367336 146946
rect 367284 146882 367336 146888
rect 368480 32428 368532 32434
rect 368480 32370 368532 32376
rect 368492 16574 368520 32370
rect 368584 18630 368612 161446
rect 368572 18624 368624 18630
rect 368572 18566 368624 18572
rect 367204 16546 367784 16574
rect 368492 16546 369440 16574
rect 367100 9308 367152 9314
rect 367100 9250 367152 9256
rect 367008 3460 367060 3466
rect 367008 3402 367060 3408
rect 367020 480 367048 3402
rect 362286 354 362398 480
rect 361868 326 362398 354
rect 362286 -960 362398 326
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 367756 354 367784 16546
rect 369412 480 369440 16546
rect 369872 4894 369900 180118
rect 370148 175658 370176 180118
rect 369964 175630 370176 175658
rect 369964 9246 369992 175630
rect 370700 161474 370728 180118
rect 370148 161446 370728 161474
rect 370148 108322 370176 161446
rect 370136 108316 370188 108322
rect 370136 108258 370188 108264
rect 370044 22840 370096 22846
rect 370044 22782 370096 22788
rect 370056 16574 370084 22782
rect 370056 16546 370176 16574
rect 369952 9240 370004 9246
rect 369952 9182 370004 9188
rect 369860 4888 369912 4894
rect 369860 4830 369912 4836
rect 368174 354 368286 480
rect 367756 326 368286 354
rect 368174 -960 368286 326
rect 369370 -960 369482 480
rect 370148 354 370176 16546
rect 371252 4826 371280 180118
rect 371620 161474 371648 180118
rect 371884 176724 371936 176730
rect 371884 176666 371936 176672
rect 371344 161446 371648 161474
rect 371344 9178 371372 161446
rect 371896 40730 371924 176666
rect 372724 175658 372752 180118
rect 372632 175630 372752 175658
rect 372816 180118 373106 180146
rect 373658 180118 373764 180146
rect 372632 106962 372660 175630
rect 372816 163538 372844 180118
rect 373736 177070 373764 180118
rect 374012 180118 374118 180146
rect 374196 180118 374670 180146
rect 374840 180118 375222 180146
rect 375576 180118 375682 180146
rect 375944 180118 376234 180146
rect 376312 180118 376694 180146
rect 376772 180118 377246 180146
rect 377324 180118 377798 180146
rect 378152 180118 378258 180146
rect 378336 180118 378810 180146
rect 378888 180118 379270 180146
rect 379624 180118 379822 180146
rect 379992 180118 380374 180146
rect 380728 180118 380834 180146
rect 381004 180118 381386 180146
rect 381464 180118 381846 180146
rect 373724 177064 373776 177070
rect 373724 177006 373776 177012
rect 374012 175624 374040 180118
rect 374012 175596 374132 175624
rect 374000 175500 374052 175506
rect 374000 175442 374052 175448
rect 372804 163532 372856 163538
rect 372804 163474 372856 163480
rect 372620 106956 372672 106962
rect 372620 106898 372672 106904
rect 372620 55888 372672 55894
rect 372620 55830 372672 55836
rect 371884 40724 371936 40730
rect 371884 40666 371936 40672
rect 372632 16574 372660 55830
rect 372632 16546 372936 16574
rect 371332 9172 371384 9178
rect 371332 9114 371384 9120
rect 371700 8968 371752 8974
rect 371700 8910 371752 8916
rect 371240 4820 371292 4826
rect 371240 4762 371292 4768
rect 371712 480 371740 8910
rect 372908 480 372936 16546
rect 374012 9110 374040 175442
rect 374104 105602 374132 175596
rect 374196 162178 374224 180118
rect 374644 177064 374696 177070
rect 374644 177006 374696 177012
rect 374184 162172 374236 162178
rect 374184 162114 374236 162120
rect 374656 130422 374684 177006
rect 374840 175506 374868 180118
rect 375380 175704 375432 175710
rect 375380 175646 375432 175652
rect 374828 175500 374880 175506
rect 374828 175442 374880 175448
rect 374644 130416 374696 130422
rect 374644 130358 374696 130364
rect 374092 105596 374144 105602
rect 374092 105538 374144 105544
rect 374092 44872 374144 44878
rect 374092 44814 374144 44820
rect 374000 9104 374052 9110
rect 374000 9046 374052 9052
rect 374104 7546 374132 44814
rect 375392 9042 375420 175646
rect 375472 175636 375524 175642
rect 375472 175578 375524 175584
rect 375484 160750 375512 175578
rect 375472 160744 375524 160750
rect 375472 160686 375524 160692
rect 375576 104174 375604 180118
rect 375944 175642 375972 180118
rect 376312 175710 376340 180118
rect 376300 175704 376352 175710
rect 376300 175646 376352 175652
rect 375932 175636 375984 175642
rect 375932 175578 375984 175584
rect 375472 104168 375524 104174
rect 375472 104110 375524 104116
rect 375564 104168 375616 104174
rect 375564 104110 375616 104116
rect 375484 16574 375512 104110
rect 376772 26926 376800 180118
rect 377324 161474 377352 180118
rect 376956 161446 377352 161474
rect 376852 127628 376904 127634
rect 376852 127570 376904 127576
rect 376760 26920 376812 26926
rect 376760 26862 376812 26868
rect 376864 16574 376892 127570
rect 376956 126274 376984 161446
rect 376944 126268 376996 126274
rect 376944 126210 376996 126216
rect 375484 16546 376064 16574
rect 376864 16546 377720 16574
rect 375380 9036 375432 9042
rect 375380 8978 375432 8984
rect 374092 7540 374144 7546
rect 374092 7482 374144 7488
rect 375288 7540 375340 7546
rect 375288 7482 375340 7488
rect 374000 5092 374052 5098
rect 374000 5034 374052 5040
rect 374012 2530 374040 5034
rect 374012 2502 374132 2530
rect 374104 480 374132 2502
rect 375300 480 375328 7482
rect 370566 354 370678 480
rect 370148 326 370678 354
rect 370566 -960 370678 326
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376036 354 376064 16546
rect 377692 480 377720 16546
rect 378152 8974 378180 180118
rect 378336 102814 378364 180118
rect 378888 161474 378916 180118
rect 379520 171760 379572 171766
rect 379520 171702 379572 171708
rect 378428 161446 378916 161474
rect 378428 159390 378456 161446
rect 378416 159384 378468 159390
rect 378416 159326 378468 159332
rect 378324 102808 378376 102814
rect 378324 102750 378376 102756
rect 379532 101454 379560 171702
rect 379624 149734 379652 180118
rect 379992 171766 380020 180118
rect 380728 176730 380756 180118
rect 380716 176724 380768 176730
rect 380716 176666 380768 176672
rect 379980 171760 380032 171766
rect 379980 171702 380032 171708
rect 380900 171760 380952 171766
rect 380900 171702 380952 171708
rect 379612 149728 379664 149734
rect 379612 149670 379664 149676
rect 379520 101448 379572 101454
rect 379520 101390 379572 101396
rect 379520 57248 379572 57254
rect 379520 57190 379572 57196
rect 378876 9376 378928 9382
rect 378876 9318 378928 9324
rect 378140 8968 378192 8974
rect 378140 8910 378192 8916
rect 378888 480 378916 9318
rect 376454 354 376566 480
rect 376036 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379532 354 379560 57190
rect 380912 44878 380940 171702
rect 381004 127634 381032 180118
rect 381464 171766 381492 180118
rect 381544 176724 381596 176730
rect 381544 176666 381596 176672
rect 381452 171760 381504 171766
rect 381452 171702 381504 171708
rect 381556 158030 381584 176666
rect 382568 176654 382596 180254
rect 382384 176626 382596 176654
rect 382660 180118 382950 180146
rect 383028 180118 383410 180146
rect 383764 180118 383962 180146
rect 384422 180118 384528 180146
rect 382384 166994 382412 176626
rect 382660 166994 382688 180118
rect 382292 166966 382412 166994
rect 382476 166966 382688 166994
rect 382292 164234 382320 166966
rect 382200 164206 382320 164234
rect 381544 158024 381596 158030
rect 381544 157966 381596 157972
rect 382200 156670 382228 164206
rect 382476 159372 382504 166966
rect 382292 159344 382504 159372
rect 382188 156664 382240 156670
rect 382188 156606 382240 156612
rect 380992 127628 381044 127634
rect 380992 127570 381044 127576
rect 380900 44872 380952 44878
rect 380900 44814 380952 44820
rect 382292 24138 382320 159344
rect 383028 157334 383056 180118
rect 383660 171692 383712 171698
rect 383660 171634 383712 171640
rect 382476 157306 383056 157334
rect 382372 60036 382424 60042
rect 382372 59978 382424 59984
rect 380900 24132 380952 24138
rect 380900 24074 380952 24080
rect 382280 24132 382332 24138
rect 382280 24074 382332 24080
rect 380912 16574 380940 24074
rect 382384 16574 382412 59978
rect 382476 42090 382504 157306
rect 383672 51746 383700 171634
rect 383764 155242 383792 180118
rect 384500 176730 384528 180118
rect 384592 180118 384974 180146
rect 385144 180118 385526 180146
rect 385696 180118 385986 180146
rect 386432 180118 386538 180146
rect 386616 180118 386998 180146
rect 387550 180118 387748 180146
rect 384488 176724 384540 176730
rect 384488 176666 384540 176672
rect 384592 171698 384620 180118
rect 385040 171760 385092 171766
rect 385040 171702 385092 171708
rect 384580 171692 384632 171698
rect 384580 171634 384632 171640
rect 383752 155236 383804 155242
rect 383752 155178 383804 155184
rect 383660 51740 383712 51746
rect 383660 51682 383712 51688
rect 382556 42220 382608 42226
rect 382556 42162 382608 42168
rect 382464 42084 382516 42090
rect 382464 42026 382516 42032
rect 380912 16546 381216 16574
rect 381188 480 381216 16546
rect 382292 16546 382412 16574
rect 382292 3466 382320 16546
rect 382568 6914 382596 42162
rect 385052 25566 385080 171702
rect 385144 153882 385172 180118
rect 385592 176724 385644 176730
rect 385592 176666 385644 176672
rect 385604 166994 385632 176666
rect 385696 171766 385724 180118
rect 385684 171760 385736 171766
rect 385684 171702 385736 171708
rect 385604 166966 385724 166994
rect 385132 153876 385184 153882
rect 385132 153818 385184 153824
rect 385696 129062 385724 166966
rect 385132 129056 385184 129062
rect 385132 128998 385184 129004
rect 385684 129056 385736 129062
rect 385684 128998 385736 129004
rect 383660 25560 383712 25566
rect 383660 25502 383712 25508
rect 385040 25560 385092 25566
rect 385040 25502 385092 25508
rect 383672 16574 383700 25502
rect 385144 16574 385172 128998
rect 386432 98666 386460 180118
rect 386616 151094 386644 180118
rect 387720 174554 387748 180118
rect 387904 180118 388102 180146
rect 388272 180118 388562 180146
rect 388732 180118 389114 180146
rect 389284 180118 389574 180146
rect 390126 180118 390416 180146
rect 387708 174548 387760 174554
rect 387708 174490 387760 174496
rect 387800 171760 387852 171766
rect 387800 171702 387852 171708
rect 386604 151088 386656 151094
rect 386604 151030 386656 151036
rect 386420 98660 386472 98666
rect 386420 98602 386472 98608
rect 386420 58676 386472 58682
rect 386420 58618 386472 58624
rect 386432 16574 386460 58618
rect 383672 16546 384344 16574
rect 385144 16546 386000 16574
rect 386432 16546 386736 16574
rect 382384 6886 382596 6914
rect 382280 3460 382332 3466
rect 382280 3402 382332 3408
rect 382384 480 382412 6886
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 383580 480 383608 3402
rect 379950 354 380062 480
rect 379532 326 380062 354
rect 379950 -960 380062 326
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384316 354 384344 16546
rect 385972 480 386000 16546
rect 384734 354 384846 480
rect 384316 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386708 354 386736 16546
rect 387812 6186 387840 171702
rect 387904 49026 387932 180118
rect 388272 171766 388300 180118
rect 388260 171760 388312 171766
rect 388260 171702 388312 171708
rect 388732 157334 388760 180118
rect 387996 157306 388760 157334
rect 387996 148374 388024 157306
rect 389180 152516 389232 152522
rect 389180 152458 389232 152464
rect 387984 148368 388036 148374
rect 387984 148310 388036 148316
rect 387892 49020 387944 49026
rect 387892 48962 387944 48968
rect 387892 26988 387944 26994
rect 387892 26930 387944 26936
rect 387800 6180 387852 6186
rect 387800 6122 387852 6128
rect 387126 354 387238 480
rect 386708 326 387238 354
rect 387904 354 387932 26930
rect 389192 16574 389220 152458
rect 389284 97306 389312 180118
rect 390388 175982 390416 180118
rect 390572 180118 390678 180146
rect 390756 180118 391138 180146
rect 391400 180118 391690 180146
rect 390376 175976 390428 175982
rect 390376 175918 390428 175924
rect 389272 97300 389324 97306
rect 389272 97242 389324 97248
rect 389192 16546 389496 16574
rect 389468 480 389496 16546
rect 390572 3194 390600 180118
rect 390652 18692 390704 18698
rect 390652 18634 390704 18640
rect 390664 3602 390692 18634
rect 390756 5234 390784 180118
rect 391400 161474 391428 180118
rect 391940 163600 391992 163606
rect 391940 163542 391992 163548
rect 390848 161446 391428 161474
rect 390744 5228 390796 5234
rect 390744 5170 390796 5176
rect 390848 3641 390876 161446
rect 391952 16574 391980 163542
rect 393320 61396 393372 61402
rect 393320 61338 393372 61344
rect 393332 16574 393360 61338
rect 393976 20670 394004 194647
rect 394068 33114 394096 204303
rect 394160 60722 394188 224975
rect 394252 73166 394280 234631
rect 394344 100706 394372 254215
rect 394436 113150 394464 264279
rect 394528 153202 394556 294335
rect 394620 193186 394648 324391
rect 395344 314764 395396 314770
rect 395344 314706 395396 314712
rect 394608 193180 394660 193186
rect 394608 193122 394660 193128
rect 394606 185056 394662 185065
rect 394606 184991 394662 185000
rect 394620 184958 394648 184991
rect 394608 184952 394660 184958
rect 394608 184894 394660 184900
rect 395356 179382 395384 314706
rect 399484 284572 399536 284578
rect 399484 284514 399536 284520
rect 396724 244588 396776 244594
rect 396724 244530 396776 244536
rect 395344 179376 395396 179382
rect 395344 179318 395396 179324
rect 394700 176044 394752 176050
rect 394700 175986 394752 175992
rect 394516 153196 394568 153202
rect 394516 153138 394568 153144
rect 394424 113144 394476 113150
rect 394424 113086 394476 113092
rect 394332 100700 394384 100706
rect 394332 100642 394384 100648
rect 394240 73160 394292 73166
rect 394240 73102 394292 73108
rect 394148 60716 394200 60722
rect 394148 60658 394200 60664
rect 394056 33108 394108 33114
rect 394056 33050 394108 33056
rect 393964 20664 394016 20670
rect 393964 20606 394016 20612
rect 394712 16574 394740 175986
rect 396080 153944 396132 153950
rect 396080 153886 396132 153892
rect 391952 16546 392624 16574
rect 393332 16546 394280 16574
rect 394712 16546 395384 16574
rect 390928 14544 390980 14550
rect 390928 14486 390980 14492
rect 390834 3632 390890 3641
rect 390652 3596 390704 3602
rect 390834 3567 390890 3576
rect 390652 3538 390704 3544
rect 390940 3482 390968 14486
rect 391020 5228 391072 5234
rect 391020 5170 391072 5176
rect 390664 3454 390968 3482
rect 391032 3466 391060 5170
rect 391848 3596 391900 3602
rect 391848 3538 391900 3544
rect 391940 3596 391992 3602
rect 391940 3538 391992 3544
rect 391020 3460 391072 3466
rect 390560 3188 390612 3194
rect 390560 3130 390612 3136
rect 390664 480 390692 3454
rect 391020 3402 391072 3408
rect 391860 480 391888 3538
rect 391952 3466 391980 3538
rect 391940 3460 391992 3466
rect 391940 3402 391992 3408
rect 392032 3460 392084 3466
rect 392032 3402 392084 3408
rect 392044 3194 392072 3402
rect 392032 3188 392084 3194
rect 392032 3130 392084 3136
rect 388230 354 388342 480
rect 387904 326 388342 354
rect 387126 -960 387238 326
rect 388230 -960 388342 326
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 392596 354 392624 16546
rect 394252 480 394280 16546
rect 395356 480 395384 16546
rect 393014 354 393126 480
rect 392596 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396092 354 396120 153886
rect 396736 86970 396764 244530
rect 398840 149796 398892 149802
rect 398840 149738 398892 149744
rect 396724 86964 396776 86970
rect 396724 86906 396776 86912
rect 397460 19984 397512 19990
rect 397460 19926 397512 19932
rect 397472 16574 397500 19926
rect 397472 16546 397776 16574
rect 397748 480 397776 16546
rect 398852 3074 398880 149738
rect 399496 139398 399524 284514
rect 406396 245614 406424 358770
rect 479536 299470 479564 361898
rect 486424 361888 486476 361894
rect 486424 361830 486476 361836
rect 483664 361820 483716 361826
rect 483664 361762 483716 361768
rect 482284 361684 482336 361690
rect 482284 361626 482336 361632
rect 482296 353258 482324 361626
rect 482284 353252 482336 353258
rect 482284 353194 482336 353200
rect 479524 299464 479576 299470
rect 479524 299406 479576 299412
rect 483676 273222 483704 361762
rect 485044 361752 485096 361758
rect 485044 361694 485096 361700
rect 485056 325650 485084 361694
rect 485044 325644 485096 325650
rect 485044 325586 485096 325592
rect 483664 273216 483716 273222
rect 483664 273158 483716 273164
rect 486436 259418 486464 361830
rect 489184 361616 489236 361622
rect 489184 361558 489236 361564
rect 489196 313274 489224 361558
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 489184 313268 489236 313274
rect 489184 313210 489236 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 554044 303680 554096 303686
rect 554044 303622 554096 303628
rect 551284 274712 551336 274718
rect 551284 274654 551336 274660
rect 486424 259412 486476 259418
rect 486424 259354 486476 259360
rect 406384 245608 406436 245614
rect 406384 245550 406436 245556
rect 457444 213988 457496 213994
rect 457444 213930 457496 213936
rect 418160 177744 418212 177750
rect 418160 177686 418212 177692
rect 407120 171896 407172 171902
rect 407120 171838 407172 171844
rect 400220 164960 400272 164966
rect 400220 164902 400272 164908
rect 399484 139392 399536 139398
rect 399484 139334 399536 139340
rect 400232 16574 400260 164902
rect 404360 155304 404412 155310
rect 404360 155246 404412 155252
rect 400232 16546 400904 16574
rect 398932 10736 398984 10742
rect 398932 10678 398984 10684
rect 398944 3194 398972 10678
rect 398932 3188 398984 3194
rect 398932 3130 398984 3136
rect 400128 3188 400180 3194
rect 400128 3130 400180 3136
rect 398852 3046 398972 3074
rect 398944 480 398972 3046
rect 400140 480 400168 3130
rect 396510 354 396622 480
rect 396092 326 396622 354
rect 396510 -960 396622 326
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 400876 354 400904 16546
rect 403624 10668 403676 10674
rect 403624 10610 403676 10616
rect 402520 6452 402572 6458
rect 402520 6394 402572 6400
rect 402532 480 402560 6394
rect 403636 480 403664 10610
rect 401294 354 401406 480
rect 400876 326 401406 354
rect 401294 -960 401406 326
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404372 354 404400 155246
rect 406016 6384 406068 6390
rect 406016 6326 406068 6332
rect 406028 480 406056 6326
rect 407132 3074 407160 171838
rect 416780 162240 416832 162246
rect 416780 162182 416832 162188
rect 411260 160812 411312 160818
rect 411260 160754 411312 160760
rect 407212 156732 407264 156738
rect 407212 156674 407264 156680
rect 407224 3194 407252 156674
rect 408500 43444 408552 43450
rect 408500 43386 408552 43392
rect 408512 16574 408540 43386
rect 411272 16574 411300 160754
rect 415492 29640 415544 29646
rect 415492 29582 415544 29588
rect 408512 16546 409184 16574
rect 411272 16546 411944 16574
rect 407212 3188 407264 3194
rect 407212 3130 407264 3136
rect 408408 3188 408460 3194
rect 408408 3130 408460 3136
rect 407132 3046 407252 3074
rect 407224 480 407252 3046
rect 408420 480 408448 3130
rect 404790 354 404902 480
rect 404372 326 404902 354
rect 404790 -960 404902 326
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409156 354 409184 16546
rect 410800 10600 410852 10606
rect 410800 10542 410852 10548
rect 410812 480 410840 10542
rect 411916 480 411944 16546
rect 414296 10532 414348 10538
rect 414296 10474 414348 10480
rect 413100 6316 413152 6322
rect 413100 6258 413152 6264
rect 413112 480 413140 6258
rect 414308 480 414336 10474
rect 415504 3262 415532 29582
rect 416792 16574 416820 162182
rect 418172 16574 418200 177686
rect 425060 177676 425112 177682
rect 425060 177618 425112 177624
rect 423680 148436 423732 148442
rect 423680 148378 423732 148384
rect 416792 16546 417464 16574
rect 418172 16546 418568 16574
rect 415400 3256 415452 3262
rect 415400 3198 415452 3204
rect 415492 3256 415544 3262
rect 415492 3198 415544 3204
rect 416688 3256 416740 3262
rect 416688 3198 416740 3204
rect 415412 1714 415440 3198
rect 415412 1686 415532 1714
rect 415504 480 415532 1686
rect 416700 480 416728 3198
rect 409574 354 409686 480
rect 409156 326 409686 354
rect 409574 -960 409686 326
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 16546
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 418540 354 418568 16546
rect 420920 10464 420972 10470
rect 420920 10406 420972 10412
rect 420184 6248 420236 6254
rect 420184 6190 420236 6196
rect 420196 480 420224 6190
rect 418958 354 419070 480
rect 418540 326 419070 354
rect 417854 -960 417966 326
rect 418958 -960 419070 326
rect 420154 -960 420266 480
rect 420932 354 420960 10406
rect 422576 3324 422628 3330
rect 422576 3266 422628 3272
rect 422588 480 422616 3266
rect 423692 3210 423720 148378
rect 425072 16574 425100 177618
rect 431960 177608 432012 177614
rect 431960 177550 432012 177556
rect 430580 147008 430632 147014
rect 430580 146950 430632 146956
rect 426440 35216 426492 35222
rect 426440 35158 426492 35164
rect 426452 16574 426480 35158
rect 430592 16574 430620 146950
rect 425072 16546 425744 16574
rect 426452 16546 426848 16574
rect 430592 16546 430896 16574
rect 423772 10396 423824 10402
rect 423772 10338 423824 10344
rect 423784 3398 423812 10338
rect 423772 3392 423824 3398
rect 423772 3334 423824 3340
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 423692 3182 423812 3210
rect 423784 480 423812 3182
rect 424980 480 425008 3334
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 425716 354 425744 16546
rect 426134 354 426246 480
rect 425716 326 426246 354
rect 426820 354 426848 16546
rect 428464 10328 428516 10334
rect 428464 10270 428516 10276
rect 428476 480 428504 10270
rect 429660 3324 429712 3330
rect 429660 3266 429712 3272
rect 429672 480 429700 3266
rect 430868 480 430896 16546
rect 431972 3398 432000 177550
rect 440240 177540 440292 177546
rect 440240 177482 440292 177488
rect 438860 159452 438912 159458
rect 438860 159394 438912 159400
rect 434720 158092 434772 158098
rect 434720 158034 434772 158040
rect 432052 124908 432104 124914
rect 432052 124850 432104 124856
rect 431960 3392 432012 3398
rect 431960 3334 432012 3340
rect 432064 480 432092 124850
rect 433340 31068 433392 31074
rect 433340 31010 433392 31016
rect 433352 16574 433380 31010
rect 434732 16574 434760 158034
rect 437480 93152 437532 93158
rect 437480 93094 437532 93100
rect 433352 16546 434024 16574
rect 434732 16546 435128 16574
rect 433248 3392 433300 3398
rect 433248 3334 433300 3340
rect 433260 480 433288 3334
rect 427238 354 427350 480
rect 426820 326 427350 354
rect 426134 -960 426246 326
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 433996 354 434024 16546
rect 434414 354 434526 480
rect 433996 326 434526 354
rect 435100 354 435128 16546
rect 436744 4140 436796 4146
rect 436744 4082 436796 4088
rect 436756 480 436784 4082
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437492 354 437520 93094
rect 438872 16574 438900 159394
rect 438872 16546 439176 16574
rect 439148 480 439176 16546
rect 440252 3210 440280 177482
rect 447140 177472 447192 177478
rect 447140 177414 447192 177420
rect 440332 145580 440384 145586
rect 440332 145522 440384 145528
rect 440344 3398 440372 145522
rect 441620 123480 441672 123486
rect 441620 123422 441672 123428
rect 441632 16574 441660 123422
rect 445760 122120 445812 122126
rect 445760 122062 445812 122068
rect 444380 28280 444432 28286
rect 444380 28222 444432 28228
rect 444392 16574 444420 28222
rect 441632 16546 442672 16574
rect 444392 16546 445064 16574
rect 440332 3392 440384 3398
rect 440332 3334 440384 3340
rect 441528 3392 441580 3398
rect 441528 3334 441580 3340
rect 440252 3182 440372 3210
rect 440344 480 440372 3182
rect 441540 480 441568 3334
rect 442644 480 442672 16546
rect 443828 4072 443880 4078
rect 443828 4014 443880 4020
rect 443840 480 443868 4014
rect 445036 480 445064 16546
rect 437910 354 438022 480
rect 437492 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 122062
rect 447152 16574 447180 177414
rect 454040 177404 454092 177410
rect 454040 177346 454092 177352
rect 448520 173256 448572 173262
rect 448520 173198 448572 173204
rect 447152 16546 447456 16574
rect 447428 480 447456 16546
rect 448532 1970 448560 173198
rect 448612 144220 448664 144226
rect 448612 144162 448664 144168
rect 448520 1964 448572 1970
rect 448520 1906 448572 1912
rect 448624 480 448652 144162
rect 452660 120760 452712 120766
rect 452660 120702 452712 120708
rect 451280 94512 451332 94518
rect 451280 94454 451332 94460
rect 451292 16574 451320 94454
rect 452672 16574 452700 120702
rect 451292 16546 451688 16574
rect 452672 16546 453344 16574
rect 450912 4004 450964 4010
rect 450912 3946 450964 3952
rect 449808 1964 449860 1970
rect 449808 1906 449860 1912
rect 449820 480 449848 1906
rect 450924 480 450952 3946
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 16546
rect 453316 480 453344 16546
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454052 354 454080 177346
rect 457456 46918 457484 213930
rect 460940 177336 460992 177342
rect 460940 177278 460992 177284
rect 459560 169108 459612 169114
rect 459560 169050 459612 169056
rect 458180 142860 458232 142866
rect 458180 142802 458232 142808
rect 457444 46912 457496 46918
rect 457444 46854 457496 46860
rect 456892 46232 456944 46238
rect 456892 46174 456944 46180
rect 455696 8016 455748 8022
rect 455696 7958 455748 7964
rect 455708 480 455736 7958
rect 456904 480 456932 46174
rect 458192 16574 458220 142802
rect 459572 16574 459600 169050
rect 460952 16574 460980 177278
rect 483020 174616 483072 174622
rect 483020 174558 483072 174564
rect 463700 119400 463752 119406
rect 463700 119342 463752 119348
rect 463712 16574 463740 119342
rect 473360 117972 473412 117978
rect 473360 117914 473412 117920
rect 458192 16546 459232 16574
rect 459572 16546 459968 16574
rect 460952 16546 461624 16574
rect 463712 16546 464016 16574
rect 458088 3936 458140 3942
rect 458088 3878 458140 3884
rect 458100 480 458128 3878
rect 459204 480 459232 16546
rect 454470 354 454582 480
rect 454052 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 16546
rect 461596 480 461624 16546
rect 462780 7948 462832 7954
rect 462780 7890 462832 7896
rect 462792 480 462820 7890
rect 463988 480 464016 16546
rect 467472 12096 467524 12102
rect 467472 12038 467524 12044
rect 466276 7880 466328 7886
rect 466276 7822 466328 7828
rect 465172 3868 465224 3874
rect 465172 3810 465224 3816
rect 465184 480 465212 3810
rect 466288 480 466316 7822
rect 467484 480 467512 12038
rect 470600 12028 470652 12034
rect 470600 11970 470652 11976
rect 469864 7812 469916 7818
rect 469864 7754 469916 7760
rect 468668 3800 468720 3806
rect 468668 3742 468720 3748
rect 468680 480 468708 3742
rect 469876 480 469904 7754
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 11970
rect 472256 3732 472308 3738
rect 472256 3674 472308 3680
rect 472268 480 472296 3674
rect 473372 3534 473400 117914
rect 481640 116612 481692 116618
rect 481640 116554 481692 116560
rect 473452 33788 473504 33794
rect 473452 33730 473504 33736
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 473464 480 473492 33730
rect 481652 16574 481680 116554
rect 483032 16574 483060 174558
rect 489920 173188 489972 173194
rect 489920 173130 489972 173136
rect 484400 141432 484452 141438
rect 484400 141374 484452 141380
rect 484412 16574 484440 141374
rect 481652 16546 482416 16574
rect 483032 16546 484072 16574
rect 484412 16546 484808 16574
rect 480536 14476 480588 14482
rect 480536 14418 480588 14424
rect 478144 11960 478196 11966
rect 478144 11902 478196 11908
rect 476948 7744 477000 7750
rect 476948 7686 477000 7692
rect 475752 3664 475804 3670
rect 475752 3606 475804 3612
rect 474188 3528 474240 3534
rect 474188 3470 474240 3476
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474200 354 474228 3470
rect 475764 480 475792 3606
rect 476960 480 476988 7686
rect 478156 480 478184 11902
rect 479340 3392 479392 3398
rect 479340 3334 479392 3340
rect 479352 480 479380 3334
rect 480548 480 480576 14418
rect 481732 7676 481784 7682
rect 481732 7618 481784 7624
rect 481744 480 481772 7618
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 16546
rect 484044 480 484072 16546
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 484780 354 484808 16546
rect 487160 15904 487212 15910
rect 487160 15846 487212 15852
rect 486424 11892 486476 11898
rect 486424 11834 486476 11840
rect 486436 480 486464 11834
rect 485198 354 485310 480
rect 484780 326 485310 354
rect 485198 -960 485310 326
rect 486394 -960 486506 480
rect 487172 354 487200 15846
rect 488816 7608 488868 7614
rect 488816 7550 488868 7556
rect 488828 480 488856 7550
rect 489932 3534 489960 173130
rect 494060 171828 494112 171834
rect 494060 171770 494112 171776
rect 490012 115252 490064 115258
rect 490012 115194 490064 115200
rect 489920 3528 489972 3534
rect 489920 3470 489972 3476
rect 490024 3346 490052 115194
rect 491300 36576 491352 36582
rect 491300 36518 491352 36524
rect 491312 16574 491340 36518
rect 494072 16574 494100 171770
rect 500960 170400 501012 170406
rect 500960 170342 501012 170348
rect 495440 140072 495492 140078
rect 495440 140014 495492 140020
rect 491312 16546 492352 16574
rect 494072 16546 494744 16574
rect 490748 3528 490800 3534
rect 490748 3470 490800 3476
rect 489932 3318 490052 3346
rect 489932 480 489960 3318
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3470
rect 492324 480 492352 16546
rect 493048 11824 493100 11830
rect 493048 11766 493100 11772
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 11766
rect 494716 480 494744 16546
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495452 354 495480 140014
rect 499580 113824 499632 113830
rect 499580 113766 499632 113772
rect 498200 22772 498252 22778
rect 498200 22714 498252 22720
rect 497096 11756 497148 11762
rect 497096 11698 497148 11704
rect 497108 480 497136 11698
rect 498212 3534 498240 22714
rect 498292 21412 498344 21418
rect 498292 21354 498344 21360
rect 498200 3528 498252 3534
rect 498200 3470 498252 3476
rect 498304 3346 498332 21354
rect 499592 16574 499620 113766
rect 500972 16574 501000 170342
rect 507860 169040 507912 169046
rect 507860 168982 507912 168988
rect 502340 137284 502392 137290
rect 502340 137226 502392 137232
rect 502352 16574 502380 137226
rect 506480 135924 506532 135930
rect 506480 135866 506532 135872
rect 505100 91792 505152 91798
rect 505100 91734 505152 91740
rect 505112 16574 505140 91734
rect 499592 16546 500632 16574
rect 500972 16546 501368 16574
rect 502352 16546 503024 16574
rect 505112 16546 505416 16574
rect 499028 3528 499080 3534
rect 499028 3470 499080 3476
rect 498212 3318 498332 3346
rect 498212 480 498240 3318
rect 495870 354 495982 480
rect 495452 326 495982 354
rect 495870 -960 495982 326
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499040 354 499068 3470
rect 500604 480 500632 16546
rect 499366 354 499478 480
rect 499040 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501340 354 501368 16546
rect 502996 480 503024 16546
rect 503720 13320 503772 13326
rect 503720 13262 503772 13268
rect 501758 354 501870 480
rect 501340 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503732 354 503760 13262
rect 505388 480 505416 16546
rect 506492 480 506520 135866
rect 506572 47592 506624 47598
rect 506572 47534 506624 47540
rect 506584 16574 506612 47534
rect 507872 16574 507900 168982
rect 514760 167680 514812 167686
rect 514760 167622 514812 167628
rect 513380 134564 513432 134570
rect 513380 134506 513432 134512
rect 509240 37936 509292 37942
rect 509240 37878 509292 37884
rect 509252 16574 509280 37878
rect 506584 16546 507256 16574
rect 507872 16546 508912 16574
rect 509252 16546 509648 16574
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 16546
rect 508884 480 508912 16546
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509620 354 509648 16546
rect 511264 13252 511316 13258
rect 511264 13194 511316 13200
rect 511276 480 511304 13194
rect 512460 5024 512512 5030
rect 512460 4966 512512 4972
rect 512472 480 512500 4966
rect 510038 354 510150 480
rect 509620 326 510150 354
rect 510038 -960 510150 326
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513392 354 513420 134506
rect 514772 3534 514800 167622
rect 525800 166320 525852 166326
rect 525800 166262 525852 166268
rect 516140 133204 516192 133210
rect 516140 133146 516192 133152
rect 514852 111104 514904 111110
rect 514852 111046 514904 111052
rect 514760 3528 514812 3534
rect 514760 3470 514812 3476
rect 514864 3346 514892 111046
rect 516152 16574 516180 133146
rect 520280 131776 520332 131782
rect 520280 131718 520332 131724
rect 516152 16546 517192 16574
rect 515588 3528 515640 3534
rect 515588 3470 515640 3476
rect 514772 3318 514892 3346
rect 514772 480 514800 3318
rect 513534 354 513646 480
rect 513392 326 513646 354
rect 513534 -960 513646 326
rect 514730 -960 514842 480
rect 515600 354 515628 3470
rect 517164 480 517192 16546
rect 517888 13184 517940 13190
rect 517888 13126 517940 13132
rect 515926 354 516038 480
rect 515600 326 516038 354
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517900 354 517928 13126
rect 519544 5024 519596 5030
rect 519544 4966 519596 4972
rect 519556 480 519584 4966
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 131718
rect 524420 109744 524472 109750
rect 524420 109686 524472 109692
rect 523040 39364 523092 39370
rect 523040 39306 523092 39312
rect 521660 13116 521712 13122
rect 521660 13058 521712 13064
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 13058
rect 523052 3534 523080 39306
rect 523132 17264 523184 17270
rect 523132 17206 523184 17212
rect 523040 3528 523092 3534
rect 523040 3470 523092 3476
rect 523144 3346 523172 17206
rect 524432 16574 524460 109686
rect 525812 16574 525840 166262
rect 529940 164892 529992 164898
rect 529940 164834 529992 164840
rect 528560 146940 528612 146946
rect 528560 146882 528612 146888
rect 524432 16546 525472 16574
rect 525812 16546 526208 16574
rect 523868 3528 523920 3534
rect 523868 3470 523920 3476
rect 523052 3318 523172 3346
rect 523052 480 523080 3318
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523880 354 523908 3470
rect 525444 480 525472 16546
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526180 354 526208 16546
rect 527824 9308 527876 9314
rect 527824 9250 527876 9256
rect 527836 480 527864 9250
rect 526598 354 526710 480
rect 526180 326 526710 354
rect 526598 -960 526710 326
rect 527794 -960 527906 480
rect 528572 354 528600 146882
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 529952 354 529980 164834
rect 539600 163532 539652 163538
rect 539600 163474 539652 163480
rect 535460 108316 535512 108322
rect 535460 108258 535512 108264
rect 531320 40724 531372 40730
rect 531320 40666 531372 40672
rect 531332 480 531360 40666
rect 531412 18624 531464 18630
rect 531412 18566 531464 18572
rect 531424 16574 531452 18566
rect 535472 16574 535500 108258
rect 531424 16546 532096 16574
rect 535472 16546 536144 16574
rect 530094 354 530206 480
rect 529952 326 530206 354
rect 528990 -960 529102 326
rect 530094 -960 530206 326
rect 531290 -960 531402 480
rect 532068 354 532096 16546
rect 534908 9240 534960 9246
rect 534908 9182 534960 9188
rect 533712 4888 533764 4894
rect 533712 4830 533764 4836
rect 533724 480 533752 4830
rect 534920 480 534948 9182
rect 536116 480 536144 16546
rect 538404 9172 538456 9178
rect 538404 9114 538456 9120
rect 537208 4820 537260 4826
rect 537208 4762 537260 4768
rect 537220 480 537248 4762
rect 538416 480 538444 9114
rect 539612 3534 539640 163474
rect 543740 162172 543792 162178
rect 543740 162114 543792 162120
rect 540980 130416 541032 130422
rect 540980 130358 541032 130364
rect 539692 106956 539744 106962
rect 539692 106898 539744 106904
rect 539600 3528 539652 3534
rect 539600 3470 539652 3476
rect 539704 3346 539732 106898
rect 540992 16574 541020 130358
rect 542360 105596 542412 105602
rect 542360 105538 542412 105544
rect 542372 16574 542400 105538
rect 543752 16574 543780 162114
rect 547880 160744 547932 160750
rect 547880 160686 547932 160692
rect 546500 104168 546552 104174
rect 546500 104110 546552 104116
rect 540992 16546 542032 16574
rect 542372 16546 542768 16574
rect 543752 16546 544424 16574
rect 540428 3528 540480 3534
rect 540428 3470 540480 3476
rect 539612 3318 539732 3346
rect 539612 480 539640 3318
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540440 354 540468 3470
rect 542004 480 542032 16546
rect 540766 354 540878 480
rect 540440 326 540878 354
rect 540766 -960 540878 326
rect 541962 -960 542074 480
rect 542740 354 542768 16546
rect 544396 480 544424 16546
rect 545488 9104 545540 9110
rect 545488 9046 545540 9052
rect 545500 480 545528 9046
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 104110
rect 547892 480 547920 160686
rect 551296 126954 551324 274654
rect 554056 167006 554084 303622
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579804 206984 579856 206990
rect 579804 206926 579856 206932
rect 579816 205737 579844 206926
rect 579802 205728 579858 205737
rect 579802 205663 579858 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 576124 184952 576176 184958
rect 576124 184894 576176 184900
rect 571984 174548 572036 174554
rect 571984 174490 572036 174496
rect 554044 167000 554096 167006
rect 554044 166942 554096 166948
rect 554780 159384 554832 159390
rect 554780 159326 554832 159332
rect 551284 126948 551336 126954
rect 551284 126890 551336 126896
rect 550640 126268 550692 126274
rect 550640 126210 550692 126216
rect 549260 26920 549312 26926
rect 549260 26862 549312 26868
rect 549272 16574 549300 26862
rect 550652 16574 550680 126210
rect 553400 102808 553452 102814
rect 553400 102750 553452 102756
rect 553412 16574 553440 102750
rect 549272 16546 550312 16574
rect 550652 16546 551048 16574
rect 553412 16546 553808 16574
rect 549076 9036 549128 9042
rect 549076 8978 549128 8984
rect 549088 480 549116 8978
rect 550284 480 550312 16546
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 16546
rect 552664 8968 552716 8974
rect 552664 8910 552716 8916
rect 552676 480 552704 8910
rect 553780 480 553808 16546
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 159326
rect 557540 158024 557592 158030
rect 557540 157966 557592 157972
rect 556160 149728 556212 149734
rect 556160 149670 556212 149676
rect 556172 480 556200 149670
rect 556252 101448 556304 101454
rect 556252 101390 556304 101396
rect 556264 16574 556292 101390
rect 557552 16574 557580 157966
rect 561680 156664 561732 156670
rect 561680 156606 561732 156612
rect 558920 127628 558972 127634
rect 558920 127570 558972 127576
rect 558932 16574 558960 127570
rect 560300 44872 560352 44878
rect 560300 44814 560352 44820
rect 560312 16574 560340 44814
rect 561692 16574 561720 156606
rect 564440 155236 564492 155242
rect 564440 155178 564492 155184
rect 563060 24132 563112 24138
rect 563060 24074 563112 24080
rect 556264 16546 556936 16574
rect 557552 16546 558592 16574
rect 558932 16546 559328 16574
rect 560312 16546 560432 16574
rect 561692 16546 562088 16574
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 556908 354 556936 16546
rect 558564 480 558592 16546
rect 557326 354 557438 480
rect 556908 326 557438 354
rect 557326 -960 557438 326
rect 558522 -960 558634 480
rect 559300 354 559328 16546
rect 559718 354 559830 480
rect 559300 326 559830 354
rect 560404 354 560432 16546
rect 562060 480 562088 16546
rect 560822 354 560934 480
rect 560404 326 560934 354
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563072 354 563100 24074
rect 564452 3534 564480 155178
rect 568580 153876 568632 153882
rect 568580 153818 568632 153824
rect 565820 129056 565872 129062
rect 565820 128998 565872 129004
rect 564532 42084 564584 42090
rect 564532 42026 564584 42032
rect 564440 3528 564492 3534
rect 564440 3470 564492 3476
rect 564544 3346 564572 42026
rect 565832 16574 565860 128998
rect 566464 51740 566516 51746
rect 566464 51682 566516 51688
rect 565832 16546 566412 16574
rect 565268 3528 565320 3534
rect 565268 3470 565320 3476
rect 566384 3482 566412 16546
rect 566476 4146 566504 51682
rect 568592 16574 568620 153818
rect 570604 98660 570656 98666
rect 570604 98602 570656 98608
rect 569960 25560 570012 25566
rect 569960 25502 570012 25508
rect 569972 16574 570000 25502
rect 568592 16546 568712 16574
rect 569972 16546 570368 16574
rect 566464 4140 566516 4146
rect 566464 4082 566516 4088
rect 568028 4140 568080 4146
rect 568028 4082 568080 4088
rect 564452 3318 564572 3346
rect 564452 480 564480 3318
rect 563214 354 563326 480
rect 563072 326 563326 354
rect 563214 -960 563326 326
rect 564410 -960 564522 480
rect 565280 354 565308 3470
rect 566384 3454 566872 3482
rect 566844 480 566872 3454
rect 568040 480 568068 4082
rect 565606 354 565718 480
rect 565280 326 565718 354
rect 565606 -960 565718 326
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 568684 354 568712 16546
rect 570340 480 570368 16546
rect 570616 3534 570644 98602
rect 570604 3528 570656 3534
rect 570604 3470 570656 3476
rect 571524 3528 571576 3534
rect 571524 3470 571576 3476
rect 571536 480 571564 3470
rect 571996 3058 572024 174490
rect 572812 151088 572864 151094
rect 572812 151030 572864 151036
rect 572824 6914 572852 151030
rect 574744 148368 574796 148374
rect 574744 148310 574796 148316
rect 574100 49020 574152 49026
rect 574100 48962 574152 48968
rect 574112 16574 574140 48962
rect 574112 16546 574692 16574
rect 572732 6886 572852 6914
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572732 480 572760 6886
rect 574664 3482 574692 16546
rect 574756 3874 574784 148310
rect 576136 6866 576164 184894
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 579620 175976 579672 175982
rect 579620 175918 579672 175924
rect 578240 97300 578292 97306
rect 578240 97242 578292 97248
rect 578252 16574 578280 97242
rect 578252 16546 578648 16574
rect 576124 6860 576176 6866
rect 576124 6802 576176 6808
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 574744 3868 574796 3874
rect 574744 3810 574796 3816
rect 574664 3454 575152 3482
rect 573916 3052 573968 3058
rect 573916 2994 573968 3000
rect 573928 480 573956 2994
rect 575124 480 575152 3454
rect 576320 480 576348 6122
rect 577412 3868 577464 3874
rect 577412 3810 577464 3816
rect 577424 480 577452 3810
rect 578620 480 578648 16546
rect 569102 354 569214 480
rect 568684 326 569214 354
rect 569102 -960 569214 326
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579632 354 579660 175918
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 579896 139392 579948 139398
rect 579894 139360 579896 139369
rect 579948 139360 579950 139369
rect 579894 139295 579950 139304
rect 579988 126948 580040 126954
rect 579988 126890 580040 126896
rect 580000 126041 580028 126890
rect 579986 126032 580042 126041
rect 579986 125967 580042 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 579894 33144 579950 33153
rect 579894 33079 579896 33088
rect 579948 33079 579950 33088
rect 579896 33050 579948 33056
rect 579896 20664 579948 20670
rect 579896 20606 579948 20612
rect 579908 19825 579936 20606
rect 579894 19816 579950 19825
rect 579894 19751 579950 19760
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 583390 3360 583446 3369
rect 583390 3295 583446 3304
rect 583404 480 583432 3295
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3330 606056 3386 606112
rect 3330 579944 3386 580000
rect 2962 527856 3018 527912
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 2870 475632 2926 475688
rect 2778 423564 2834 423600
rect 2778 423544 2780 423564
rect 2780 423544 2832 423564
rect 2832 423544 2834 423564
rect 3330 410488 3386 410544
rect 3330 371320 3386 371376
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3606 566888 3662 566944
rect 3698 553832 3754 553888
rect 3790 501744 3846 501800
rect 3882 462576 3938 462632
rect 3974 449520 4030 449576
rect 4066 397432 4122 397488
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 2778 319232 2834 319288
rect 3054 293120 3110 293176
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 2778 214920 2834 214976
rect 3054 201864 3110 201920
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 149776 3386 149832
rect 3054 136720 3110 136776
rect 3330 110608 3386 110664
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 2870 32408 2926 32464
rect 3606 97552 3662 97608
rect 189722 354728 189778 354784
rect 189078 344256 189134 344312
rect 189078 334328 189134 334384
rect 189078 324400 189134 324456
rect 189078 304272 189134 304328
rect 189078 274760 189134 274816
rect 189078 254224 189134 254280
rect 189078 244316 189134 244352
rect 189078 244296 189080 244316
rect 189080 244296 189132 244316
rect 189132 244296 189134 244316
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 394146 354728 394202 354784
rect 394054 344256 394110 344312
rect 393962 334328 394018 334384
rect 190090 314744 190146 314800
rect 189998 294344 190054 294400
rect 189906 264288 189962 264344
rect 189814 234640 189870 234696
rect 189078 225004 189134 225040
rect 189078 224984 189080 225004
rect 189080 224984 189132 225004
rect 189132 224984 189134 225004
rect 189078 214240 189134 214296
rect 189722 204312 189778 204368
rect 189078 194656 189134 194712
rect 3514 58520 3570 58576
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 138846 3304 138902 3360
rect 190182 284280 190238 284336
rect 190090 185000 190146 185056
rect 393778 244588 393834 244624
rect 393778 244568 393780 244588
rect 393780 244568 393832 244588
rect 393832 244568 393834 244588
rect 394606 324400 394662 324456
rect 394330 314764 394386 314800
rect 394330 314744 394332 314764
rect 394332 314744 394384 314764
rect 394384 314744 394386 314764
rect 394330 304272 394386 304328
rect 394514 294344 394570 294400
rect 394422 284572 394478 284608
rect 394422 284552 394424 284572
rect 394424 284552 394476 284572
rect 394476 284552 394478 284572
rect 394422 274760 394478 274816
rect 394422 264288 394478 264344
rect 394330 254224 394386 254280
rect 394238 234640 394294 234696
rect 394146 224984 394202 225040
rect 394054 214376 394110 214432
rect 394054 204312 394110 204368
rect 393962 194656 394018 194712
rect 197358 3304 197414 3360
rect 394606 185000 394662 185056
rect 390834 3576 390890 3632
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 579802 205672 579858 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 579894 139340 579896 139360
rect 579896 139340 579948 139360
rect 579948 139340 579950 139360
rect 579894 139304 579950 139340
rect 579986 125976 580042 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 579894 33108 579950 33144
rect 579894 33088 579896 33108
rect 579896 33088 579948 33108
rect 579948 33088 579950 33108
rect 579894 19760 579950 19816
rect 580170 6568 580226 6624
rect 583390 3304 583446 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3325 606114 3391 606117
rect -960 606112 3391 606114
rect -960 606056 3330 606112
rect 3386 606056 3391 606112
rect -960 606054 3391 606056
rect -960 605964 480 606054
rect 3325 606051 3391 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3601 566946 3667 566949
rect -960 566944 3667 566946
rect -960 566888 3606 566944
rect 3662 566888 3667 566944
rect -960 566886 3667 566888
rect -960 566796 480 566886
rect 3601 566883 3667 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3785 501802 3851 501805
rect -960 501800 3851 501802
rect -960 501744 3790 501800
rect 3846 501744 3851 501800
rect -960 501742 3851 501744
rect -960 501652 480 501742
rect 3785 501739 3851 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2865 475690 2931 475693
rect -960 475688 2931 475690
rect -960 475632 2870 475688
rect 2926 475632 2931 475688
rect -960 475630 2931 475632
rect -960 475540 480 475630
rect 2865 475627 2931 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3877 462634 3943 462637
rect -960 462632 3943 462634
rect -960 462576 3882 462632
rect 3938 462576 3943 462632
rect -960 462574 3943 462576
rect -960 462484 480 462574
rect 3877 462571 3943 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3969 449578 4035 449581
rect -960 449576 4035 449578
rect -960 449520 3974 449576
rect 4030 449520 4035 449576
rect -960 449518 4035 449520
rect -960 449428 480 449518
rect 3969 449515 4035 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 4061 397490 4127 397493
rect -960 397488 4127 397490
rect -960 397432 4066 397488
rect 4122 397432 4127 397488
rect -960 397430 4127 397432
rect -960 397340 480 397430
rect 4061 397427 4127 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 189717 354786 189783 354789
rect 192158 354786 192218 354960
rect 189717 354784 192218 354786
rect 189717 354728 189722 354784
rect 189778 354728 192218 354784
rect 189717 354726 192218 354728
rect 391798 354786 391858 354960
rect 394141 354786 394207 354789
rect 391798 354784 394207 354786
rect 391798 354728 394146 354784
rect 394202 354728 394207 354784
rect 391798 354726 394207 354728
rect 189717 354723 189783 354726
rect 394141 354723 394207 354726
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 189073 344314 189139 344317
rect 192158 344314 192218 344896
rect 189073 344312 192218 344314
rect 189073 344256 189078 344312
rect 189134 344256 192218 344312
rect 189073 344254 192218 344256
rect 391798 344314 391858 344896
rect 394049 344314 394115 344317
rect 391798 344312 394115 344314
rect 391798 344256 394054 344312
rect 394110 344256 394115 344312
rect 391798 344254 394115 344256
rect 189073 344251 189139 344254
rect 394049 344251 394115 344254
rect 583520 338452 584960 338692
rect 189073 334386 189139 334389
rect 192158 334386 192218 334968
rect 189073 334384 192218 334386
rect 189073 334328 189078 334384
rect 189134 334328 192218 334384
rect 189073 334326 192218 334328
rect 391798 334386 391858 334968
rect 393957 334386 394023 334389
rect 391798 334384 394023 334386
rect 391798 334328 393962 334384
rect 394018 334328 394023 334384
rect 391798 334326 394023 334328
rect 189073 334323 189139 334326
rect 393957 334323 394023 334326
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 189073 324458 189139 324461
rect 192158 324458 192218 324904
rect 189073 324456 192218 324458
rect 189073 324400 189078 324456
rect 189134 324400 192218 324456
rect 189073 324398 192218 324400
rect 391798 324458 391858 324904
rect 394601 324458 394667 324461
rect 391798 324456 394667 324458
rect 391798 324400 394606 324456
rect 394662 324400 394667 324456
rect 391798 324398 394667 324400
rect 189073 324395 189139 324398
rect 394601 324395 394667 324398
rect -960 319290 480 319380
rect 2773 319290 2839 319293
rect -960 319288 2839 319290
rect -960 319232 2778 319288
rect 2834 319232 2839 319288
rect -960 319230 2839 319232
rect -960 319140 480 319230
rect 2773 319227 2839 319230
rect 190085 314802 190151 314805
rect 192158 314802 192218 314976
rect 190085 314800 192218 314802
rect 190085 314744 190090 314800
rect 190146 314744 192218 314800
rect 190085 314742 192218 314744
rect 391798 314802 391858 314976
rect 394325 314802 394391 314805
rect 391798 314800 394391 314802
rect 391798 314744 394330 314800
rect 394386 314744 394391 314800
rect 391798 314742 394391 314744
rect 190085 314739 190151 314742
rect 394325 314739 394391 314742
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 189073 304330 189139 304333
rect 192158 304330 192218 304912
rect 189073 304328 192218 304330
rect 189073 304272 189078 304328
rect 189134 304272 192218 304328
rect 189073 304270 192218 304272
rect 391798 304330 391858 304912
rect 394325 304330 394391 304333
rect 391798 304328 394391 304330
rect 391798 304272 394330 304328
rect 394386 304272 394391 304328
rect 391798 304270 394391 304272
rect 189073 304267 189139 304270
rect 394325 304267 394391 304270
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 189993 294402 190059 294405
rect 192158 294402 192218 294984
rect 189993 294400 192218 294402
rect 189993 294344 189998 294400
rect 190054 294344 192218 294400
rect 189993 294342 192218 294344
rect 391798 294402 391858 294984
rect 394509 294402 394575 294405
rect 391798 294400 394575 294402
rect 391798 294344 394514 294400
rect 394570 294344 394575 294400
rect 391798 294342 394575 294344
rect 189993 294339 190059 294342
rect 394509 294339 394575 294342
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 583520 285276 584960 285516
rect 190177 284338 190243 284341
rect 192158 284338 192218 284920
rect 391798 284610 391858 284920
rect 394417 284610 394483 284613
rect 391798 284608 394483 284610
rect 391798 284552 394422 284608
rect 394478 284552 394483 284608
rect 391798 284550 394483 284552
rect 394417 284547 394483 284550
rect 190177 284336 192218 284338
rect 190177 284280 190182 284336
rect 190238 284280 192218 284336
rect 190177 284278 192218 284280
rect 190177 284275 190243 284278
rect -960 279972 480 280212
rect 189073 274818 189139 274821
rect 192158 274818 192218 274992
rect 189073 274816 192218 274818
rect 189073 274760 189078 274816
rect 189134 274760 192218 274816
rect 189073 274758 192218 274760
rect 391798 274818 391858 274992
rect 394417 274818 394483 274821
rect 391798 274816 394483 274818
rect 391798 274760 394422 274816
rect 394478 274760 394483 274816
rect 391798 274758 394483 274760
rect 189073 274755 189139 274758
rect 394417 274755 394483 274758
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 189901 264346 189967 264349
rect 192158 264346 192218 264928
rect 189901 264344 192218 264346
rect 189901 264288 189906 264344
rect 189962 264288 192218 264344
rect 189901 264286 192218 264288
rect 391798 264346 391858 264928
rect 394417 264346 394483 264349
rect 391798 264344 394483 264346
rect 391798 264288 394422 264344
rect 394478 264288 394483 264344
rect 391798 264286 394483 264288
rect 189901 264283 189967 264286
rect 394417 264283 394483 264286
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 189073 254282 189139 254285
rect 192158 254282 192218 254864
rect 189073 254280 192218 254282
rect -960 254146 480 254236
rect 189073 254224 189078 254280
rect 189134 254224 192218 254280
rect 189073 254222 192218 254224
rect 391798 254282 391858 254864
rect 394325 254282 394391 254285
rect 391798 254280 394391 254282
rect 391798 254224 394330 254280
rect 394386 254224 394391 254280
rect 391798 254222 394391 254224
rect 189073 254219 189139 254222
rect 394325 254219 394391 254222
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 189073 244354 189139 244357
rect 192158 244354 192218 244936
rect 391798 244626 391858 244936
rect 393773 244626 393839 244629
rect 391798 244624 393839 244626
rect 391798 244568 393778 244624
rect 393834 244568 393839 244624
rect 391798 244566 393839 244568
rect 393773 244563 393839 244566
rect 189073 244352 192218 244354
rect 189073 244296 189078 244352
rect 189134 244296 192218 244352
rect 189073 244294 192218 244296
rect 189073 244291 189139 244294
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 189809 234698 189875 234701
rect 192158 234698 192218 234872
rect 189809 234696 192218 234698
rect 189809 234640 189814 234696
rect 189870 234640 192218 234696
rect 189809 234638 192218 234640
rect 391798 234698 391858 234872
rect 394233 234698 394299 234701
rect 391798 234696 394299 234698
rect 391798 234640 394238 234696
rect 394294 234640 394299 234696
rect 391798 234638 394299 234640
rect 189809 234635 189875 234638
rect 394233 234635 394299 234638
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 189073 225042 189139 225045
rect 394141 225042 394207 225045
rect 189073 225040 192218 225042
rect 189073 224984 189078 225040
rect 189134 224984 192218 225040
rect 189073 224982 192218 224984
rect 189073 224979 189139 224982
rect 192158 224944 192218 224982
rect 391798 225040 394207 225042
rect 391798 224984 394146 225040
rect 394202 224984 394207 225040
rect 391798 224982 394207 224984
rect 391798 224944 391858 224982
rect 394141 224979 394207 224982
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 189073 214298 189139 214301
rect 192158 214298 192218 214880
rect 391798 214434 391858 214880
rect 394049 214434 394115 214437
rect 391798 214432 394115 214434
rect 391798 214376 394054 214432
rect 394110 214376 394115 214432
rect 391798 214374 394115 214376
rect 394049 214371 394115 214374
rect 189073 214296 192218 214298
rect 189073 214240 189078 214296
rect 189134 214240 192218 214296
rect 189073 214238 192218 214240
rect 189073 214235 189139 214238
rect 579797 205730 579863 205733
rect 583520 205730 584960 205820
rect 579797 205728 584960 205730
rect 579797 205672 579802 205728
rect 579858 205672 584960 205728
rect 579797 205670 584960 205672
rect 579797 205667 579863 205670
rect 583520 205580 584960 205670
rect 189717 204370 189783 204373
rect 192158 204370 192218 204952
rect 189717 204368 192218 204370
rect 189717 204312 189722 204368
rect 189778 204312 192218 204368
rect 189717 204310 192218 204312
rect 391798 204370 391858 204952
rect 394049 204370 394115 204373
rect 391798 204368 394115 204370
rect 391798 204312 394054 204368
rect 394110 204312 394115 204368
rect 391798 204310 394115 204312
rect 189717 204307 189783 204310
rect 394049 204307 394115 204310
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 189073 194714 189139 194717
rect 192158 194714 192218 194888
rect 189073 194712 192218 194714
rect 189073 194656 189078 194712
rect 189134 194656 192218 194712
rect 189073 194654 192218 194656
rect 391798 194714 391858 194888
rect 393957 194714 394023 194717
rect 391798 194712 394023 194714
rect 391798 194656 393962 194712
rect 394018 194656 394023 194712
rect 391798 194654 394023 194656
rect 189073 194651 189139 194654
rect 393957 194651 394023 194654
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 190085 185058 190151 185061
rect 394601 185058 394667 185061
rect 190085 185056 192218 185058
rect 190085 185000 190090 185056
rect 190146 185000 192218 185056
rect 190085 184998 192218 185000
rect 190085 184995 190151 184998
rect 192158 184960 192218 184998
rect 391798 185056 394667 185058
rect 391798 185000 394606 185056
rect 394662 185000 394667 185056
rect 391798 184998 394667 185000
rect 391798 184960 391858 184998
rect 394601 184995 394667 184998
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3325 149834 3391 149837
rect -960 149832 3391 149834
rect -960 149776 3330 149832
rect 3386 149776 3391 149832
rect -960 149774 3391 149776
rect -960 149684 480 149774
rect 3325 149771 3391 149774
rect 579889 139362 579955 139365
rect 583520 139362 584960 139452
rect 579889 139360 584960 139362
rect 579889 139304 579894 139360
rect 579950 139304 584960 139360
rect 579889 139302 584960 139304
rect 579889 139299 579955 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 579981 126034 580047 126037
rect 583520 126034 584960 126124
rect 579981 126032 584960 126034
rect 579981 125976 579986 126032
rect 580042 125976 584960 126032
rect 579981 125974 584960 125976
rect 579981 125971 580047 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 579889 33146 579955 33149
rect 583520 33146 584960 33236
rect 579889 33144 584960 33146
rect 579889 33088 579894 33144
rect 579950 33088 584960 33144
rect 579889 33086 584960 33088
rect 579889 33083 579955 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 579889 19818 579955 19821
rect 583520 19818 584960 19908
rect 579889 19816 584960 19818
rect 579889 19760 579894 19816
rect 579950 19760 584960 19816
rect 579889 19758 584960 19760
rect 579889 19755 579955 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 390829 3634 390895 3637
rect 390829 3632 393330 3634
rect 390829 3576 390834 3632
rect 390890 3576 393330 3632
rect 390829 3574 393330 3576
rect 390829 3571 390895 3574
rect 138841 3362 138907 3365
rect 197353 3362 197419 3365
rect 138841 3360 197419 3362
rect 138841 3304 138846 3360
rect 138902 3304 197358 3360
rect 197414 3304 197419 3360
rect 138841 3302 197419 3304
rect 393270 3362 393330 3574
rect 583385 3362 583451 3365
rect 393270 3360 583451 3362
rect 393270 3304 583390 3360
rect 583446 3304 583451 3360
rect 393270 3302 583451 3304
rect 138841 3299 138907 3302
rect 197353 3299 197419 3302
rect 583385 3299 583451 3302
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 381454 92414 416898
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 385174 96134 420618
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 362000 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 362000 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 362000 204134 384618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 362000 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 362000 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 362000 218414 362898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 362000 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 362000 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 362000 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 362000 236414 380898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 362000 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 362000 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 362000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 362000 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 362000 258134 366618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 362000 261854 370338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 362000 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 362000 272414 380898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 362000 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 362000 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 362000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 362000 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 362000 294134 366618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 362000 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 362000 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 362000 308414 380898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 362000 312134 384618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 362000 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 362000 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 362000 326414 362898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 362000 330134 366618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 362000 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 362000 337574 374058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 362000 344414 380898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 362000 348134 384618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 362000 351854 388338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 362000 355574 392058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 362000 362414 362898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 362000 366134 366618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 362000 369854 370338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 362000 373574 374058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 362000 380414 380898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 362000 384134 384618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 362000 387854 388338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 362000 391574 392058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 211568 345454 211888 345486
rect 211568 345218 211610 345454
rect 211846 345218 211888 345454
rect 211568 345134 211888 345218
rect 211568 344898 211610 345134
rect 211846 344898 211888 345134
rect 211568 344866 211888 344898
rect 242288 345454 242608 345486
rect 242288 345218 242330 345454
rect 242566 345218 242608 345454
rect 242288 345134 242608 345218
rect 242288 344898 242330 345134
rect 242566 344898 242608 345134
rect 242288 344866 242608 344898
rect 273008 345454 273328 345486
rect 273008 345218 273050 345454
rect 273286 345218 273328 345454
rect 273008 345134 273328 345218
rect 273008 344898 273050 345134
rect 273286 344898 273328 345134
rect 273008 344866 273328 344898
rect 303728 345454 304048 345486
rect 303728 345218 303770 345454
rect 304006 345218 304048 345454
rect 303728 345134 304048 345218
rect 303728 344898 303770 345134
rect 304006 344898 304048 345134
rect 303728 344866 304048 344898
rect 334448 345454 334768 345486
rect 334448 345218 334490 345454
rect 334726 345218 334768 345454
rect 334448 345134 334768 345218
rect 334448 344898 334490 345134
rect 334726 344898 334768 345134
rect 334448 344866 334768 344898
rect 365168 345454 365488 345486
rect 365168 345218 365210 345454
rect 365446 345218 365488 345454
rect 365168 345134 365488 345218
rect 365168 344898 365210 345134
rect 365446 344898 365488 345134
rect 365168 344866 365488 344898
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 196208 327454 196528 327486
rect 196208 327218 196250 327454
rect 196486 327218 196528 327454
rect 196208 327134 196528 327218
rect 196208 326898 196250 327134
rect 196486 326898 196528 327134
rect 196208 326866 196528 326898
rect 226928 327454 227248 327486
rect 226928 327218 226970 327454
rect 227206 327218 227248 327454
rect 226928 327134 227248 327218
rect 226928 326898 226970 327134
rect 227206 326898 227248 327134
rect 226928 326866 227248 326898
rect 257648 327454 257968 327486
rect 257648 327218 257690 327454
rect 257926 327218 257968 327454
rect 257648 327134 257968 327218
rect 257648 326898 257690 327134
rect 257926 326898 257968 327134
rect 257648 326866 257968 326898
rect 288368 327454 288688 327486
rect 288368 327218 288410 327454
rect 288646 327218 288688 327454
rect 288368 327134 288688 327218
rect 288368 326898 288410 327134
rect 288646 326898 288688 327134
rect 288368 326866 288688 326898
rect 319088 327454 319408 327486
rect 319088 327218 319130 327454
rect 319366 327218 319408 327454
rect 319088 327134 319408 327218
rect 319088 326898 319130 327134
rect 319366 326898 319408 327134
rect 319088 326866 319408 326898
rect 349808 327454 350128 327486
rect 349808 327218 349850 327454
rect 350086 327218 350128 327454
rect 349808 327134 350128 327218
rect 349808 326898 349850 327134
rect 350086 326898 350128 327134
rect 349808 326866 350128 326898
rect 380528 327454 380848 327486
rect 380528 327218 380570 327454
rect 380806 327218 380848 327454
rect 380528 327134 380848 327218
rect 380528 326898 380570 327134
rect 380806 326898 380848 327134
rect 380528 326866 380848 326898
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 211568 309454 211888 309486
rect 211568 309218 211610 309454
rect 211846 309218 211888 309454
rect 211568 309134 211888 309218
rect 211568 308898 211610 309134
rect 211846 308898 211888 309134
rect 211568 308866 211888 308898
rect 242288 309454 242608 309486
rect 242288 309218 242330 309454
rect 242566 309218 242608 309454
rect 242288 309134 242608 309218
rect 242288 308898 242330 309134
rect 242566 308898 242608 309134
rect 242288 308866 242608 308898
rect 273008 309454 273328 309486
rect 273008 309218 273050 309454
rect 273286 309218 273328 309454
rect 273008 309134 273328 309218
rect 273008 308898 273050 309134
rect 273286 308898 273328 309134
rect 273008 308866 273328 308898
rect 303728 309454 304048 309486
rect 303728 309218 303770 309454
rect 304006 309218 304048 309454
rect 303728 309134 304048 309218
rect 303728 308898 303770 309134
rect 304006 308898 304048 309134
rect 303728 308866 304048 308898
rect 334448 309454 334768 309486
rect 334448 309218 334490 309454
rect 334726 309218 334768 309454
rect 334448 309134 334768 309218
rect 334448 308898 334490 309134
rect 334726 308898 334768 309134
rect 334448 308866 334768 308898
rect 365168 309454 365488 309486
rect 365168 309218 365210 309454
rect 365446 309218 365488 309454
rect 365168 309134 365488 309218
rect 365168 308898 365210 309134
rect 365446 308898 365488 309134
rect 365168 308866 365488 308898
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 196208 291454 196528 291486
rect 196208 291218 196250 291454
rect 196486 291218 196528 291454
rect 196208 291134 196528 291218
rect 196208 290898 196250 291134
rect 196486 290898 196528 291134
rect 196208 290866 196528 290898
rect 226928 291454 227248 291486
rect 226928 291218 226970 291454
rect 227206 291218 227248 291454
rect 226928 291134 227248 291218
rect 226928 290898 226970 291134
rect 227206 290898 227248 291134
rect 226928 290866 227248 290898
rect 257648 291454 257968 291486
rect 257648 291218 257690 291454
rect 257926 291218 257968 291454
rect 257648 291134 257968 291218
rect 257648 290898 257690 291134
rect 257926 290898 257968 291134
rect 257648 290866 257968 290898
rect 288368 291454 288688 291486
rect 288368 291218 288410 291454
rect 288646 291218 288688 291454
rect 288368 291134 288688 291218
rect 288368 290898 288410 291134
rect 288646 290898 288688 291134
rect 288368 290866 288688 290898
rect 319088 291454 319408 291486
rect 319088 291218 319130 291454
rect 319366 291218 319408 291454
rect 319088 291134 319408 291218
rect 319088 290898 319130 291134
rect 319366 290898 319408 291134
rect 319088 290866 319408 290898
rect 349808 291454 350128 291486
rect 349808 291218 349850 291454
rect 350086 291218 350128 291454
rect 349808 291134 350128 291218
rect 349808 290898 349850 291134
rect 350086 290898 350128 291134
rect 349808 290866 350128 290898
rect 380528 291454 380848 291486
rect 380528 291218 380570 291454
rect 380806 291218 380848 291454
rect 380528 291134 380848 291218
rect 380528 290898 380570 291134
rect 380806 290898 380848 291134
rect 380528 290866 380848 290898
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 211568 273454 211888 273486
rect 211568 273218 211610 273454
rect 211846 273218 211888 273454
rect 211568 273134 211888 273218
rect 211568 272898 211610 273134
rect 211846 272898 211888 273134
rect 211568 272866 211888 272898
rect 242288 273454 242608 273486
rect 242288 273218 242330 273454
rect 242566 273218 242608 273454
rect 242288 273134 242608 273218
rect 242288 272898 242330 273134
rect 242566 272898 242608 273134
rect 242288 272866 242608 272898
rect 273008 273454 273328 273486
rect 273008 273218 273050 273454
rect 273286 273218 273328 273454
rect 273008 273134 273328 273218
rect 273008 272898 273050 273134
rect 273286 272898 273328 273134
rect 273008 272866 273328 272898
rect 303728 273454 304048 273486
rect 303728 273218 303770 273454
rect 304006 273218 304048 273454
rect 303728 273134 304048 273218
rect 303728 272898 303770 273134
rect 304006 272898 304048 273134
rect 303728 272866 304048 272898
rect 334448 273454 334768 273486
rect 334448 273218 334490 273454
rect 334726 273218 334768 273454
rect 334448 273134 334768 273218
rect 334448 272898 334490 273134
rect 334726 272898 334768 273134
rect 334448 272866 334768 272898
rect 365168 273454 365488 273486
rect 365168 273218 365210 273454
rect 365446 273218 365488 273454
rect 365168 273134 365488 273218
rect 365168 272898 365210 273134
rect 365446 272898 365488 273134
rect 365168 272866 365488 272898
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 196208 255454 196528 255486
rect 196208 255218 196250 255454
rect 196486 255218 196528 255454
rect 196208 255134 196528 255218
rect 196208 254898 196250 255134
rect 196486 254898 196528 255134
rect 196208 254866 196528 254898
rect 226928 255454 227248 255486
rect 226928 255218 226970 255454
rect 227206 255218 227248 255454
rect 226928 255134 227248 255218
rect 226928 254898 226970 255134
rect 227206 254898 227248 255134
rect 226928 254866 227248 254898
rect 257648 255454 257968 255486
rect 257648 255218 257690 255454
rect 257926 255218 257968 255454
rect 257648 255134 257968 255218
rect 257648 254898 257690 255134
rect 257926 254898 257968 255134
rect 257648 254866 257968 254898
rect 288368 255454 288688 255486
rect 288368 255218 288410 255454
rect 288646 255218 288688 255454
rect 288368 255134 288688 255218
rect 288368 254898 288410 255134
rect 288646 254898 288688 255134
rect 288368 254866 288688 254898
rect 319088 255454 319408 255486
rect 319088 255218 319130 255454
rect 319366 255218 319408 255454
rect 319088 255134 319408 255218
rect 319088 254898 319130 255134
rect 319366 254898 319408 255134
rect 319088 254866 319408 254898
rect 349808 255454 350128 255486
rect 349808 255218 349850 255454
rect 350086 255218 350128 255454
rect 349808 255134 350128 255218
rect 349808 254898 349850 255134
rect 350086 254898 350128 255134
rect 349808 254866 350128 254898
rect 380528 255454 380848 255486
rect 380528 255218 380570 255454
rect 380806 255218 380848 255454
rect 380528 255134 380848 255218
rect 380528 254898 380570 255134
rect 380806 254898 380848 255134
rect 380528 254866 380848 254898
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 211568 237454 211888 237486
rect 211568 237218 211610 237454
rect 211846 237218 211888 237454
rect 211568 237134 211888 237218
rect 211568 236898 211610 237134
rect 211846 236898 211888 237134
rect 211568 236866 211888 236898
rect 242288 237454 242608 237486
rect 242288 237218 242330 237454
rect 242566 237218 242608 237454
rect 242288 237134 242608 237218
rect 242288 236898 242330 237134
rect 242566 236898 242608 237134
rect 242288 236866 242608 236898
rect 273008 237454 273328 237486
rect 273008 237218 273050 237454
rect 273286 237218 273328 237454
rect 273008 237134 273328 237218
rect 273008 236898 273050 237134
rect 273286 236898 273328 237134
rect 273008 236866 273328 236898
rect 303728 237454 304048 237486
rect 303728 237218 303770 237454
rect 304006 237218 304048 237454
rect 303728 237134 304048 237218
rect 303728 236898 303770 237134
rect 304006 236898 304048 237134
rect 303728 236866 304048 236898
rect 334448 237454 334768 237486
rect 334448 237218 334490 237454
rect 334726 237218 334768 237454
rect 334448 237134 334768 237218
rect 334448 236898 334490 237134
rect 334726 236898 334768 237134
rect 334448 236866 334768 236898
rect 365168 237454 365488 237486
rect 365168 237218 365210 237454
rect 365446 237218 365488 237454
rect 365168 237134 365488 237218
rect 365168 236898 365210 237134
rect 365446 236898 365488 237134
rect 365168 236866 365488 236898
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 196208 219454 196528 219486
rect 196208 219218 196250 219454
rect 196486 219218 196528 219454
rect 196208 219134 196528 219218
rect 196208 218898 196250 219134
rect 196486 218898 196528 219134
rect 196208 218866 196528 218898
rect 226928 219454 227248 219486
rect 226928 219218 226970 219454
rect 227206 219218 227248 219454
rect 226928 219134 227248 219218
rect 226928 218898 226970 219134
rect 227206 218898 227248 219134
rect 226928 218866 227248 218898
rect 257648 219454 257968 219486
rect 257648 219218 257690 219454
rect 257926 219218 257968 219454
rect 257648 219134 257968 219218
rect 257648 218898 257690 219134
rect 257926 218898 257968 219134
rect 257648 218866 257968 218898
rect 288368 219454 288688 219486
rect 288368 219218 288410 219454
rect 288646 219218 288688 219454
rect 288368 219134 288688 219218
rect 288368 218898 288410 219134
rect 288646 218898 288688 219134
rect 288368 218866 288688 218898
rect 319088 219454 319408 219486
rect 319088 219218 319130 219454
rect 319366 219218 319408 219454
rect 319088 219134 319408 219218
rect 319088 218898 319130 219134
rect 319366 218898 319408 219134
rect 319088 218866 319408 218898
rect 349808 219454 350128 219486
rect 349808 219218 349850 219454
rect 350086 219218 350128 219454
rect 349808 219134 350128 219218
rect 349808 218898 349850 219134
rect 350086 218898 350128 219134
rect 349808 218866 350128 218898
rect 380528 219454 380848 219486
rect 380528 219218 380570 219454
rect 380806 219218 380848 219454
rect 380528 219134 380848 219218
rect 380528 218898 380570 219134
rect 380806 218898 380848 219134
rect 380528 218866 380848 218898
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 211568 201454 211888 201486
rect 211568 201218 211610 201454
rect 211846 201218 211888 201454
rect 211568 201134 211888 201218
rect 211568 200898 211610 201134
rect 211846 200898 211888 201134
rect 211568 200866 211888 200898
rect 242288 201454 242608 201486
rect 242288 201218 242330 201454
rect 242566 201218 242608 201454
rect 242288 201134 242608 201218
rect 242288 200898 242330 201134
rect 242566 200898 242608 201134
rect 242288 200866 242608 200898
rect 273008 201454 273328 201486
rect 273008 201218 273050 201454
rect 273286 201218 273328 201454
rect 273008 201134 273328 201218
rect 273008 200898 273050 201134
rect 273286 200898 273328 201134
rect 273008 200866 273328 200898
rect 303728 201454 304048 201486
rect 303728 201218 303770 201454
rect 304006 201218 304048 201454
rect 303728 201134 304048 201218
rect 303728 200898 303770 201134
rect 304006 200898 304048 201134
rect 303728 200866 304048 200898
rect 334448 201454 334768 201486
rect 334448 201218 334490 201454
rect 334726 201218 334768 201454
rect 334448 201134 334768 201218
rect 334448 200898 334490 201134
rect 334726 200898 334768 201134
rect 334448 200866 334768 200898
rect 365168 201454 365488 201486
rect 365168 201218 365210 201454
rect 365446 201218 365488 201454
rect 365168 201134 365488 201218
rect 365168 200898 365210 201134
rect 365446 200898 365488 201134
rect 365168 200866 365488 200898
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 196208 183454 196528 183486
rect 196208 183218 196250 183454
rect 196486 183218 196528 183454
rect 196208 183134 196528 183218
rect 196208 182898 196250 183134
rect 196486 182898 196528 183134
rect 196208 182866 196528 182898
rect 226928 183454 227248 183486
rect 226928 183218 226970 183454
rect 227206 183218 227248 183454
rect 226928 183134 227248 183218
rect 226928 182898 226970 183134
rect 227206 182898 227248 183134
rect 226928 182866 227248 182898
rect 257648 183454 257968 183486
rect 257648 183218 257690 183454
rect 257926 183218 257968 183454
rect 257648 183134 257968 183218
rect 257648 182898 257690 183134
rect 257926 182898 257968 183134
rect 257648 182866 257968 182898
rect 288368 183454 288688 183486
rect 288368 183218 288410 183454
rect 288646 183218 288688 183454
rect 288368 183134 288688 183218
rect 288368 182898 288410 183134
rect 288646 182898 288688 183134
rect 288368 182866 288688 182898
rect 319088 183454 319408 183486
rect 319088 183218 319130 183454
rect 319366 183218 319408 183454
rect 319088 183134 319408 183218
rect 319088 182898 319130 183134
rect 319366 182898 319408 183134
rect 319088 182866 319408 182898
rect 349808 183454 350128 183486
rect 349808 183218 349850 183454
rect 350086 183218 350128 183454
rect 349808 183134 350128 183218
rect 349808 182898 349850 183134
rect 350086 182898 350128 183134
rect 349808 182866 350128 182898
rect 380528 183454 380848 183486
rect 380528 183218 380570 183454
rect 380806 183218 380848 183454
rect 380528 183134 380848 183218
rect 380528 182898 380570 183134
rect 380806 182898 380848 183134
rect 380528 182866 380848 182898
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 158614 193574 178000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 165454 200414 178000
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 169174 204134 178000
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 172894 207854 178000
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 178000
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 147454 218414 178000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 151174 222134 178000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 154894 225854 178000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 158614 229574 178000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 165454 236414 178000
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 169174 240134 178000
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 178000
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 178000
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 178000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 151174 258134 178000
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 154894 261854 178000
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 178000
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 165454 272414 178000
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 178000
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 178000
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 176614 283574 178000
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 147454 290414 178000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 151174 294134 178000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 154894 297854 178000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 158614 301574 178000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 165454 308414 178000
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 178000
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 178000
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 178000
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 147454 326414 178000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 151174 330134 178000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 154894 333854 178000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 158614 337574 178000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 165454 344414 178000
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 169174 348134 178000
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 172894 351854 178000
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 176614 355574 178000
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 147454 362414 178000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 151174 366134 178000
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 154894 369854 178000
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 158614 373574 178000
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 165454 380414 178000
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 169174 384134 178000
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 172894 387854 178000
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 176614 391574 178000
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 211610 345218 211846 345454
rect 211610 344898 211846 345134
rect 242330 345218 242566 345454
rect 242330 344898 242566 345134
rect 273050 345218 273286 345454
rect 273050 344898 273286 345134
rect 303770 345218 304006 345454
rect 303770 344898 304006 345134
rect 334490 345218 334726 345454
rect 334490 344898 334726 345134
rect 365210 345218 365446 345454
rect 365210 344898 365446 345134
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 196250 327218 196486 327454
rect 196250 326898 196486 327134
rect 226970 327218 227206 327454
rect 226970 326898 227206 327134
rect 257690 327218 257926 327454
rect 257690 326898 257926 327134
rect 288410 327218 288646 327454
rect 288410 326898 288646 327134
rect 319130 327218 319366 327454
rect 319130 326898 319366 327134
rect 349850 327218 350086 327454
rect 349850 326898 350086 327134
rect 380570 327218 380806 327454
rect 380570 326898 380806 327134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 211610 309218 211846 309454
rect 211610 308898 211846 309134
rect 242330 309218 242566 309454
rect 242330 308898 242566 309134
rect 273050 309218 273286 309454
rect 273050 308898 273286 309134
rect 303770 309218 304006 309454
rect 303770 308898 304006 309134
rect 334490 309218 334726 309454
rect 334490 308898 334726 309134
rect 365210 309218 365446 309454
rect 365210 308898 365446 309134
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 196250 291218 196486 291454
rect 196250 290898 196486 291134
rect 226970 291218 227206 291454
rect 226970 290898 227206 291134
rect 257690 291218 257926 291454
rect 257690 290898 257926 291134
rect 288410 291218 288646 291454
rect 288410 290898 288646 291134
rect 319130 291218 319366 291454
rect 319130 290898 319366 291134
rect 349850 291218 350086 291454
rect 349850 290898 350086 291134
rect 380570 291218 380806 291454
rect 380570 290898 380806 291134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 211610 273218 211846 273454
rect 211610 272898 211846 273134
rect 242330 273218 242566 273454
rect 242330 272898 242566 273134
rect 273050 273218 273286 273454
rect 273050 272898 273286 273134
rect 303770 273218 304006 273454
rect 303770 272898 304006 273134
rect 334490 273218 334726 273454
rect 334490 272898 334726 273134
rect 365210 273218 365446 273454
rect 365210 272898 365446 273134
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 196250 255218 196486 255454
rect 196250 254898 196486 255134
rect 226970 255218 227206 255454
rect 226970 254898 227206 255134
rect 257690 255218 257926 255454
rect 257690 254898 257926 255134
rect 288410 255218 288646 255454
rect 288410 254898 288646 255134
rect 319130 255218 319366 255454
rect 319130 254898 319366 255134
rect 349850 255218 350086 255454
rect 349850 254898 350086 255134
rect 380570 255218 380806 255454
rect 380570 254898 380806 255134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 211610 237218 211846 237454
rect 211610 236898 211846 237134
rect 242330 237218 242566 237454
rect 242330 236898 242566 237134
rect 273050 237218 273286 237454
rect 273050 236898 273286 237134
rect 303770 237218 304006 237454
rect 303770 236898 304006 237134
rect 334490 237218 334726 237454
rect 334490 236898 334726 237134
rect 365210 237218 365446 237454
rect 365210 236898 365446 237134
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 196250 219218 196486 219454
rect 196250 218898 196486 219134
rect 226970 219218 227206 219454
rect 226970 218898 227206 219134
rect 257690 219218 257926 219454
rect 257690 218898 257926 219134
rect 288410 219218 288646 219454
rect 288410 218898 288646 219134
rect 319130 219218 319366 219454
rect 319130 218898 319366 219134
rect 349850 219218 350086 219454
rect 349850 218898 350086 219134
rect 380570 219218 380806 219454
rect 380570 218898 380806 219134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 211610 201218 211846 201454
rect 211610 200898 211846 201134
rect 242330 201218 242566 201454
rect 242330 200898 242566 201134
rect 273050 201218 273286 201454
rect 273050 200898 273286 201134
rect 303770 201218 304006 201454
rect 303770 200898 304006 201134
rect 334490 201218 334726 201454
rect 334490 200898 334726 201134
rect 365210 201218 365446 201454
rect 365210 200898 365446 201134
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 196250 183218 196486 183454
rect 196250 182898 196486 183134
rect 226970 183218 227206 183454
rect 226970 182898 227206 183134
rect 257690 183218 257926 183454
rect 257690 182898 257926 183134
rect 288410 183218 288646 183454
rect 288410 182898 288646 183134
rect 319130 183218 319366 183454
rect 319130 182898 319366 183134
rect 349850 183218 350086 183454
rect 349850 182898 350086 183134
rect 380570 183218 380806 183454
rect 380570 182898 380806 183134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 211610 345454
rect 211846 345218 242330 345454
rect 242566 345218 273050 345454
rect 273286 345218 303770 345454
rect 304006 345218 334490 345454
rect 334726 345218 365210 345454
rect 365446 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 211610 345134
rect 211846 344898 242330 345134
rect 242566 344898 273050 345134
rect 273286 344898 303770 345134
rect 304006 344898 334490 345134
rect 334726 344898 365210 345134
rect 365446 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 196250 327454
rect 196486 327218 226970 327454
rect 227206 327218 257690 327454
rect 257926 327218 288410 327454
rect 288646 327218 319130 327454
rect 319366 327218 349850 327454
rect 350086 327218 380570 327454
rect 380806 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 196250 327134
rect 196486 326898 226970 327134
rect 227206 326898 257690 327134
rect 257926 326898 288410 327134
rect 288646 326898 319130 327134
rect 319366 326898 349850 327134
rect 350086 326898 380570 327134
rect 380806 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 211610 309454
rect 211846 309218 242330 309454
rect 242566 309218 273050 309454
rect 273286 309218 303770 309454
rect 304006 309218 334490 309454
rect 334726 309218 365210 309454
rect 365446 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 211610 309134
rect 211846 308898 242330 309134
rect 242566 308898 273050 309134
rect 273286 308898 303770 309134
rect 304006 308898 334490 309134
rect 334726 308898 365210 309134
rect 365446 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 196250 291454
rect 196486 291218 226970 291454
rect 227206 291218 257690 291454
rect 257926 291218 288410 291454
rect 288646 291218 319130 291454
rect 319366 291218 349850 291454
rect 350086 291218 380570 291454
rect 380806 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 196250 291134
rect 196486 290898 226970 291134
rect 227206 290898 257690 291134
rect 257926 290898 288410 291134
rect 288646 290898 319130 291134
rect 319366 290898 349850 291134
rect 350086 290898 380570 291134
rect 380806 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 211610 273454
rect 211846 273218 242330 273454
rect 242566 273218 273050 273454
rect 273286 273218 303770 273454
rect 304006 273218 334490 273454
rect 334726 273218 365210 273454
rect 365446 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 211610 273134
rect 211846 272898 242330 273134
rect 242566 272898 273050 273134
rect 273286 272898 303770 273134
rect 304006 272898 334490 273134
rect 334726 272898 365210 273134
rect 365446 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 196250 255454
rect 196486 255218 226970 255454
rect 227206 255218 257690 255454
rect 257926 255218 288410 255454
rect 288646 255218 319130 255454
rect 319366 255218 349850 255454
rect 350086 255218 380570 255454
rect 380806 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 196250 255134
rect 196486 254898 226970 255134
rect 227206 254898 257690 255134
rect 257926 254898 288410 255134
rect 288646 254898 319130 255134
rect 319366 254898 349850 255134
rect 350086 254898 380570 255134
rect 380806 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 211610 237454
rect 211846 237218 242330 237454
rect 242566 237218 273050 237454
rect 273286 237218 303770 237454
rect 304006 237218 334490 237454
rect 334726 237218 365210 237454
rect 365446 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 211610 237134
rect 211846 236898 242330 237134
rect 242566 236898 273050 237134
rect 273286 236898 303770 237134
rect 304006 236898 334490 237134
rect 334726 236898 365210 237134
rect 365446 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 196250 219454
rect 196486 219218 226970 219454
rect 227206 219218 257690 219454
rect 257926 219218 288410 219454
rect 288646 219218 319130 219454
rect 319366 219218 349850 219454
rect 350086 219218 380570 219454
rect 380806 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 196250 219134
rect 196486 218898 226970 219134
rect 227206 218898 257690 219134
rect 257926 218898 288410 219134
rect 288646 218898 319130 219134
rect 319366 218898 349850 219134
rect 350086 218898 380570 219134
rect 380806 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 211610 201454
rect 211846 201218 242330 201454
rect 242566 201218 273050 201454
rect 273286 201218 303770 201454
rect 304006 201218 334490 201454
rect 334726 201218 365210 201454
rect 365446 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 211610 201134
rect 211846 200898 242330 201134
rect 242566 200898 273050 201134
rect 273286 200898 303770 201134
rect 304006 200898 334490 201134
rect 334726 200898 365210 201134
rect 365446 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 196250 183454
rect 196486 183218 226970 183454
rect 227206 183218 257690 183454
rect 257926 183218 288410 183454
rect 288646 183218 319130 183454
rect 319366 183218 349850 183454
rect 350086 183218 380570 183454
rect 380806 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 196250 183134
rect 196486 182898 226970 183134
rect 227206 182898 257690 183134
rect 257926 182898 288410 183134
rect 288646 182898 319130 183134
rect 319366 182898 349850 183134
rect 350086 182898 380570 183134
rect 380806 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use actuator_driver_controller  mprj
timestamp 0
transform 1 0 192000 0 1 180000
box 0 0 200000 180000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 362000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 362000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 362000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 362000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 362000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 362000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 362000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 362000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 362000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 362000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 362000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 362000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 362000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 362000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 362000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 362000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 362000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 362000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 362000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 362000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 362000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 362000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 362000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 362000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 362000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 362000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 362000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 362000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 362000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 362000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 362000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 362000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 362000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 362000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 362000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 362000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 362000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 362000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 362000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 362000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 362000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 362000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 362000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 362000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 362000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
