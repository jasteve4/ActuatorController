// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * spi_mod
 *
 *
 *-------------------------------------------------------------
 */
module sync_n(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif
  input wire signal_n,
  output wire signal_sn,
  input wire clock
);
  reg [3:0] signal_state;

  always@(posedge clock)
  begin
    if(signal_n)
    begin
      signal_state <= 3'b111;
    end
    else
    begin
      signal_state <= {signal_state[2:0],signal_n};
    end
  end

  assign signal_sn = signal_state == 3'b000 ? 1'b0:1'b1;


endmodule
